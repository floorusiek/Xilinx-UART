`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "W-2024.09-SP1 -- Dec 03, 2024"
`protect key_keyowner = "Xilinx"
`protect key_keyname = "xilinxt_2023_11"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
gximP30K58XOxSmZD5pmqmeyWGOrOp4Qb2WjBylngEiCq78G+ER3Tcre5kKgtkrt
WYAK99xVpllBMhiyt3y1Tt3mSB82+6ihQBi5iJERv2SfYGWlfxvw6cbf+GbWY4/i
T94DSVGjdQCXvXBfUN0KrDrN3FX13wOl//G/QdRQYrq6Ow8VX0+h5YH8QAQvlN9r
VF6pqymUIF1XWNAGHIWAqRpaEpuk75LjiIiSoizsPC814we/KXq7rem7YOMpIy0q
AgEXqTYiC6iDRhvIZDgeD0X6QkmG2dPOOb/bj3uiOPFchmtfxpv43DWZV+V5DCCf
kqKlKg2eha/M1Jv7+vf/XQ==
`protect key_keyowner = "Siemens"
`protect key_keyname = "SIEMENS-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
ZL104PRiPQ/FY2qJSrxZbvGkZAXIfm/UoUEmyfmlOoEFGUT/njgnA/vFjUCmgsmq
DmjKxn50MBPmeD+A3QYKAz4+9SG8uhuWVY7xqZoxjvUUE3sZeOUsbFcFU5yGWOgi
XJiZXuO4UO/p8dhnYnnQBXd84bcqJwmKImUcUTqJ7j+ZqpxtYvoyv8CnByfs+nhk
brb4borMIdIbpq/kTKT1e56G/iCc8mWDP7sUqQZ07gj2Lyg7rQsd4HFc8J/wa3ZM
9XAbb+z316D8umZkizdxABS9edclaRXszwe+q4RIfP/LXBdbhTLNocaF5kpDqaRz
+si352/Uy7JyMU9/REtCIA==
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ZxHSUSNR8qh4GkAJh4dlF9tMB/KOCHTUmZCQuLfZk3wJvk3HXhUl0PLzHjCXbge1
R7UKOjL1JprIHIYTMv9QaregD8brgTnpp/FQX5eAOMPz7JVIcSQ6jc6OIAf1AvgV
Xs+t+solVBlr7tMj0gGeO/2ZM7jiX+pPeWM2YnpyHaU=
`protect data_method = "aes256-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 138272)
`protect data_block
bowr/EUi2r7ByKLBYzRJEutGZCtWhFu2ziDprexaTqY012tJWY2CWobOljXNWGZq
2qcZLNd6Hn/jnZogyL1DsWbqWOPOyEWpPpafb52pspX7ZTdfcL2HqI/TAOIkDAvh
7O6a7h5ChsI1ZJ0nYOVqA5oD+VMv3jJLyMrt7QxsHliCDnWY2NVqfU8vAoZA1jh5
UngdWEwXDy94JcJFr3k7btsxkPAlMsIu1Lq0ozCRK0FyRkEaLP5HtZxWV0N5dCYW
FcfTZFoz/n7Lwn6SwTw6C8XI47NtGwmq31ikeCJdiI1NIfjOdM3Qkj2X2KSdTf7z
l7yxAZA93xH9tJ6Orj/Hl6YnjuSUJuyzo+tB5w2ikBrR7nw/3KcW5PjEISHPixNR
AStfEAatOTkg5yciK9ujwYU6YYyCuOJk9dxloSLSxrlHXnpbmTYpI7af0EiiKQmh
zo6CN86gR4Xb6eZNfdGQa+el7SO5HRg7JOVZyygeaaAPCcKHVfVHHdH+yrHeLiW7
mGv5MUJnAxIKhh0cFbE5TckFF9kntM+8xHq7vo5s2XNiLvP/2hZtxM/LHDcXl2rS
q2RJ20USH1Ms7ph4fJ0rkUw+IBb75pNA90MF6KBBNd8W0dSkhTrWr1CLjgxLDDQC
DSlcfZz+ikyYb3gcz3PYuE7hmyJzIaq3UDH1sh4PjpnKW1bP2Ps8H+VyKa52wKjk
BFnteUN7+9Sh4m9i9F9OJlXw50gepC2h7WnTYS9LAsd/GXBbZbO3yhAA1HT1tQ6j
pSg06ZY6l6TYw1AyPxRkzBbT5vC7ZonabZyJTxkUj3Efz5Rgbar7hU/YLfXGzEmd
RUEmgIqr93vkXJrZkHFDWcPkekXLd3ayaScbKuvUe5m34kXW5XHgWcx313952P95
7tl658tQojh79AmVluw9hk9fz+L5/qPnfdTsiMIAX2nYKIO4/UVkUwdK67t6jbBD
pkIFAbz2vzDCNaUvURWQyXyZ8trXgG8i4CnfxZhbMnUMsn8zOEjYWKjVoKSkIh4K
Jneb3EOI5PAR8fJxoK/1pIq4MqxaTvqkntFslL3ImmjggQtqkQ0NbMH84ud2fRmf
yGkq6PjFWl1uvEqfHmvwS7oAFtBIBcLcx0Zy0PGQg+t9BpT0fa8aHGNVHKthSucs
PW8TBYLl8R5oet2MWxCA2hEfjWTwuITjn2xuB4hNAwwxJAZwJjYQUPYiW3kiHqnL
iVe9XT1w3q96oS/6CpqUhzC2T1rj/590yCovMxANAzG8u6bhw+8cYZ4MFC0DCnli
fPqESAYi/F5qCYuilojaCcGp9Hl0Ye59TrpMUhmQsgRrE5uF+r/BHesDHhzJPCVE
mVZQSO22fdgzz4yg9inj5Xm0Ib412NLT6tYR1xo8pFDcC+IIXP0voHJkA0NgVVow
pYut5SmNm7gogZk9thrcs+z40JWgQhxs/48DAqzywkzBJPv1JC+kHhc/JOcWGZVJ
YqE3hM+swayg9aeUhtdxec9UV0tK1hUHyzjerjePcY7s0I5YF6zwoBpzPNatkvDk
wZjLSm9EDAeeouMQPIM58YMDS0clODVYmAsC1VD0bNdEJhvPI3mxBkiMdIXiC7y2
YVuu0/Dq8zLzOxfJXzQNfFJeYHo9wTHFBDArrET4DEK0Sq7BTaGGoKwea5X6ZjEu
Hdy6nub5EK1/uVLTRb34aYbF64ez/yRG/AKa0I99jCgtsNEna2vLb9H94cELNxks
YqLUr4F+PH7jahqktLeMd0JiSMX9Aob2Aeq01kNE8+1XzXlY7l/FZqtGkb5u3sOS
LrVxnkpm5o2DUvVo+6/GTLPMwxmJTsEp9GV0eL6pS/pcFtIgyEofdyh/HXoYMsYN
QwK14btmnEDYX0HRWhzIk/6OUngZWU7EgHrdCSKV+0pX8/Hzd4o961Qq3h3FlTY6
D78CLnYNhS2G/oJN+jGSS9Pcc7DQFrmq/44YGstSurQ/4W42uV9WUmenzjczvm5p
F6Z8R6drYU5dc8O9nmz0JckswZwG6VvR8QPsrVs9NrSujRLLMd2+vDoBQz+9Jq0G
Y/fzChm8eftnfKmflHagCrskwi/1JgfgO0wbPao/4i1zrE+XJ6VzYFV11QTSds75
o7X8LfYuSKpQIPoRb2FEzIKosElQikibgFTUNbweNr1iZSh3naoYDwQV8uYxIk6g
EIrLU2g7qtz5lzC4d4i6KBx0b4X4meZW4q3L283C9zlhDnwz76DTYeEP1V9pddS2
Q81rQrK2OkiFuzR2yA/K3jwEN1mhT5i1gCCULzMGbHjbz92zHYnTK3lFZ9+42Px/
G4Hz2E48zJInG/PXOGec3QbAi9w8Hiy6kq/PjoRusPxbzbK3ZJ3SKF8x4eppEJ2O
T3joPCXdTBXrxlcXqRp4uZ7PC4p54+I3qA2n/KJGh1GJvMg5dsciXBf/7c3TgkmY
TFrP15zHrNHyPgj03sF1d//rYZcCn+vxxxoUTnVQInF7yOPX09+6Rgpm2/+C5gBi
rl+HLMzddJP54lIDLJ1gsQHasQYdCL0V/JkRFS5md+z3vgnpgUmFU4YwQjYJZnUk
PqZLrgpZsAsVP3av823JXFWFaspH2iJKeq51E/ZBZCsa3TrSI+fjwd52Ule+KR6/
HUuzWTCVaCX7YEGY571vtIgCTt3svMsWLzoZIdA5SDZfv0qd4ocYHpXC2HzrDYIt
mn5CXy8f7r4jqrA2kyJRgqb/+VwxxlE6ISd222MNOswAwv9vMmx7JpJenmRMMu2w
b+zSaD74bQbuP0nJ6ynVV9VQMlpzgA1h8+zN2gfxgXYemRe+LEAtWiy8Ig0c288i
5bDVMqve7QXA9WYE1IATCCYcT8p6Wx9sK8JT5FNz6FekJnbb2AOTgxrHARkhiggV
XcG1kNg+OzAOr4gJkBic5EdCnrxHeciXHqDU1jeycmDiHEUXk2Jt23BjceI1fsaP
rGKIdsbpnHWMDqL+B87iTT7fP+nGSagnPl4+6yjilqn8w1JEj8Hl5Gocp/3QHnN8
sYCirNZEijB0SxdV1eQTR228vpZakBdOdK6yXVZ5e5XK+l1CnQwLIuqF+67RxDjV
0VbOggm+QnrnPFME56sudYuHaVPhR1URCfWLSse20brIVWSYd4GqwhZbZ7JSG43s
aPkVao4DVKAyUs2jDazT+F4T8J6/ej5mtEJSxaScuTPotroYOiRAgbDxazh9oHDu
dCqWhYUZYBozVybbPIFxEDIyqLZ1Gad5Y2AH9YiXctPXdlvKcz33Sx0ZR1U9vzFc
8esCHC/81tpB7lV2xtgfwF73Z5EFRGiEKyQt5cDPSs8ybeZuOdEuTiPCHESA8TKd
adbS62FfQe5Qe/YSL4IwoJoK6mxK5NFhp9dpRECK7MP5u33jdXgJpkWlbQIKo0cf
oJ2qZrRDZoM4YjF19e4pDKp9VkjBOvxv8CoTQHAYo0FuHa6ORAtFYIT/W3NF7kDw
RYx4jsLZqR9gwKakyyD044e4Wf5MD5U8Es/kUErdB+nytKxeYqO6XjAa7rtmaPgD
FXbc0lXEPPQzj/E8zDjXSLDEq8OiEzXL710AIsMF8pVmjRFBF6z1uANN8vgm3wlX
ntWMR8imNvJ72/KKaSHrHtC/ZFw4U7Yw1nQYNOHHCyYA3DWoWQCKyfnZZ84HxQzL
koKPVj6xL6+FreaWBQHi4WP0z5TwYeUXMSEiIBfmIXt5qu5x4kBQ765vhMfsSeK1
BaYlu4CXHUaGeC+aBGU5dS4Gf4o3a99M1OtC34fSOu2K3g4l47ARu36f7qjYU+6k
EXL4RydDNsAMSfwNiEuQYoNmYx5KIz40/Pjcg7KW9tsvGjnu+DtaOfpvbfg6N6n8
cZsRZnQhr74jwXrhxCuiAdxd/o3BKzyhX/Om2KwhIOoYWcthJMbwcS8uovkJUycc
xcJeTTmT1SCWMjpdG+mKxQXIgejA73NperAdu4nJTA2LGGHTS3V822Ki+x02L3Jj
iUPXVbV+yPdVAa7uCs2uvmUsz6yLnFWAIezuVlB6CojDOvwXQBz/1S37y8ZUuVuR
PlvwmCXGNbtradVJojEUQ1WeW/9FZmx3FwO5nGtBOckuKoc9PrFPpE+pB5qen+uz
pWs+xaq9+Sh38AFW870nvy1UiNOMnvt+2diIiIXXzZz/I8APguxdhUTlog0LWUuO
c08ALw5fVM5LV5IDvFQ7uTySkqLPnxqw+sCvhRVM4/YIyplaM8d1ssyfcgwUW7mc
tSghNF0sjx3r5dB06B6CHD//4GbD2YkYSNlJ7zkebEVJI0VlDdVuo+AJiRJxZ6G9
q3/iDqEuzf4uCHiTvrlwcscv1xATH8k5Aylu0y7FPtY2t6c9oSkegqQGDjZtwIem
bAt9xdUZb9eEMha+64IyIHF7fJWPlUMIQUffVxp/xotzzXWFT/xuSy68OgW3O+C3
HYpasu91g23WYYry4pzWWeS6smiqUwPGmCbKqc+4NE7uCII3DAmNriIlveY/iFaI
XLuiCfKceeMIHPTTffZGLKnlvUJQaSJflPXB1ebUiwFmx4S1yBvllThsmEfAT6wL
mu5W7pxe6wRsjCpgPecQ4tu+sVs54QtY0phknUJ7uiJ6ygCGB5en3upBG/ksvZLB
N9j3v+l2njgcqTCVM/SMnzyAPBMz1NX7nXU/oPGW6PQWq7JPBA/MVnhqGzWJLOQ0
SJBMyMwFzUOxLZxoydUh2anTtC58DA+kH1zSIUnrwJMydorUTqpOeQtZ5h9VOk3+
1X+rMq4l8w+6X97uoBN+OTrkUeSYacKg1rRaFJNRrn8pVS9t2ReDAyrD1oqC8nhF
FixlM8nxIma38Z7SDvry6o0QEYTx0L8Un0asO9mgVNOhg5UojXHj2du8s7KGyncw
S5ufuICbyg/UNzZYU1jP62XM1nPCsTehH63QtBRtH41xk9RH4/orHANYrP0sZUyw
vqQ9edNqkH/vEBNMgkyzGbfTi3iwqzm3CO8qgHpV6oVw4R0Ieg4tmTDFXO1T1KSS
Jf+mK8Y/a4VlhrQads2ofKoH0OqM18asNj6u/1Ncm9t3cAA+zhAACA6OILe/5sPd
B8HpPZjSStbjRtmKRZ+upXdKxlNUCFmXqzsfjm64qFULKoc0aaKtTxCKUB9kGvS5
1nXx7KqgPqbgxK328jh4lipFuS3laMRIsAgPF2xT9NGaor0SetNDmjUPCQa54mEG
eURNO0CYmFL36IbT9nR/bIK4y2TdHKC5a0M74TVr+UrQbsM1BvJVFvlvgqrJvP07
prqqMrVZ6z/8Z7DpEodBLoyqcdQhL7HTnCN9g0m0i1JSgWqObOeGlsBokBuA/C9q
n23x062EdFbqar67M6PNN8Yby6V9xb1AN4XBT855IQhGelVSwv73o+Kq9mL6JhXH
vjrHLg1sTeyF0VSVZRKGkFeQXH2rEW2dV3qpx24R+Bz+4xFHTu1dCT1EOTttP53N
ngi2022Iu4aSfCki0WGzLJ71lnXqdGQHxvhmSFG2lONev8mur0/Q4z3gFhm4tWPs
jE0P25GJwhXZ0f0bq1LCqE/2EYPspayijncjCHiSfN5lr/UeDigCO09M2EqTap4K
wiupqsVIlkAqlaKXI2mWFqhek1PTsPbT7qLLxAYOHLMJ/Rc2obVY/Xgru546rGI2
c6N2QXmo0ur0cZBJzEBvYniPVvduqxmtGaGMAH42v5shXanlx9rfzS6SElnUdmYu
Gyr9yevuk+LCitd0HDbbXGjVEyioBtRuz0worJI8wW15EQknwfugYXhamQ4hXGBr
pOQbJoyx6Qtzb6P+fiWDJ/nyTEvwbmZCVKgX2NOg02IxLMHo/Gt25N+rJ228SXsE
mXf/IUzdkmClicE0vTBvVXMh7dKWkqxmOKOHQKqz7AtrXR+UwGquaQbhswU9V/1h
MQU3y2nN9Yd0oqzIsgsHUsBiTowIV9XMLlYf4rS86JhqTTro/epkfiA7va4elsQX
yN4mxSSLv8oR8ovqpTCNugGbb4j0/OjdCCYLDSxQBoYbcTsFZZ5KGyZODH+XDXtj
YMgACEjk9iKDRFuOtEKWcGeRvf3YRe9BwyReSGGan68nXxPUMFmeffgTwN7qWEgs
M1X2hlzpjqv4k/ghDBsGLByH15rX/3X0c41uVuv7xhsNb/vJKA7d0jGc+Sa3/7Rv
UuqPv2ySHvla259Zr0+gCHfaFdZFxmGrzAMtU2b7MpvofDzCt9Ji3von/qxtbg9Z
1keb6Qds6KbwnAaLKarvS4i9MH8Zn7D7jEBxqDdFh0cskoomH41hbPbyGKkOyf46
xz15LmJSdWDxwcwstEthr+IChV4jRmN6TVL+z7rD70k2Jg2oItpTaOVAz9S81r59
eBUhjDtHo802/6jeCaq/ch+QQOgEC3TdrwAP+QWnc1IgjD25+aPjQOl90fZzQMUe
fOpkxTWqNPKSdrj7o4xs2UwSpENFB/tNxq9UjTEYeqnlrt7XwdLYeEhUkDOiTeVX
qMtF4K+9LapwPe/l+kOd8IDqlKiKRimHSnczEBpAnNdORV8pLkIEV8Femj6TvM7Y
3uQOSESiX7kS5EKewNLnNb/n++zfH4JzxsEwgdsmv/b7XPK14w3rt68xXg2GsnbW
lrv+rQfYhMLK8BtbYqnt9DVeHOeQg03BIhIT7s/M7RtYziigi9qspJ8fpJv8YrNu
wke4iUvS+7fgYp8xkZnKFFQ2TAYHotOtHdxULgoJXoLH7RnNvOS7glN9nM8Tt60/
ofxcR0/PnWolyz+mkh8D0EVy98zyYbXlUmvz059BoX91KElrmWEr5lndxzpG7TnI
4els0De03t0uW4fGZHKJ2m+QYH1nCwgvSOBpXZhC7f3y6inaxbY86JWisfKIWWHD
8k0IMh8QjBkiwiaC8Y2ZOQcm9Zj0SAeeuRbNzs1TlDZ3lAhUnoViTC4BmFXCAzp3
VyYUnQhuURi9mDPy60+3ECuAXWg7WDSeyZqRGPyn/knw3kQB2rxu+WrEsltRURez
7vJmzGiLchfzFpR2dzK0K5lFKbQwHwOjREuYYogpCMup5i0GuD2kufD59PH/HOy+
yArvONQSDdSQeD/LOuXXXwDHxF/ifnYPmt6vh849/Wvwv6jvLSrLr2Dkbr/ArDFN
0Tl4sPsw0SWuYaUvfEOaR7vHmyEa48wP2Im5umsRQUZ7aYjbwsj/0xcFtZBNrxt2
lmAXV7DFhHvn+My5bCGUxYerlq4/UILRBaHh5WKNOU1O2tTWmzYX9mfHzRvc8F/w
Fhb6jXn3MJRv87uPRID4/k9qM0H+e5FHyDkWUN9TI2C3phjT5cAUoGDWErdutWVE
x7lJ4ywRZoy/Gvv9L5EUoACGUsZVd4vipqrwXm4g0yzQ6/fvQSuNio6AKmUQ02fF
VruudThcs/YNfgPktMTrT/7PQ0PNudkFDONAu+V37EeRL9F9TtMBaW0d6/hSCsij
qJmiYi6P3hN3ot+Q3h2ZAdrH4t7toJFklAGdMMym0s5iA0mZQEkB/VqTZx8bmrCP
gCwn89YlmmNfYpjKQKm7m8Bv5VdX95sc549MUaglR8Efe4u7h4g+KyhLbulasvBo
YknMKVgSubwur+H1wVie7bJ4SMmK9+tTZcLdLJjLNr4z60U9r8JEGnADwot7Kg3M
WYmNg0hdLA1uvgQ9Uu1Hg+LYA3hGZDRFWb9ZaTAa6G18BNSJIeUcb6GcTyN6iiMf
oBiKdB3nGcKbMErtyCh7M3JLdAlxo4E2U8Y/MZdmTWLNrdXIalC8dzlaD2hzN/zl
yluZdFpcwG25suqQR5ICRl517zEaHryruEQvYWJ0bt5JiQy7ntbtbWWQZzAaTj8Q
6iCOncljlFMjLflk1tSyzRJuv+b3kCJ4mMF196+Ipd0zyHMPsPYoBsPS5kVhtwQ3
wLPj1EYSQk0n5ktAXizm5zzWH8UPzFD6A2Xm/cdWFkpc3Fbbxy/Lq+C6wWVcyOVq
UMYLJBl+WVCBxTma5JarGZrhhliZQnpIhPZ237mf041SdgS0VV53imUNeCSxOp3t
55TFUIKnGEPzPRAxS2Ug9vjMY89NpJKMs/U9nqmU/caElAJaBJC3fMB27WcwuLxG
UniiqFvavFMBvd1a6bTtikP3cRuZcb9bAdx4N5BjT1NeVEtXayCNgNGHGihMOa30
XWnKXDsAOPb8haeYt12CQwEvxYp30356zvCcOhy9XdfAgkT8Sks/DdfZGWoXGKJK
3Iqm9CCQSdpH2LGxn82U8rmPPCrCS7yHWR4gFdIB0M5DzUHOIrva1mbte6JlwC8C
nFkAp1Es5PewevjdV9N8mhxnnYwEWi5XpJkHlSxYsx2bjHjz3PorR4+g88TGn+G8
KF7uQPmpiZjDe/K2iRPq2t4jmjTCGiVW+dhvCg2rD4lgqfgiD+IynOBv968Obm4i
+wUDyTObK25rdMDcmlbTszV0pfbmUukjRl6GgSYkFiV1GH+9KCSA7qVvOfCgbbdr
E8uF+GtSCbhLPqC9JsPnguE8oTVqhpupeYQLtLOE/vP0JG06gIgEW2o6IJkXv3G0
OJN7t/rWV4QwBSTBiUBw29XkLrU+Y5XORq4/k/ljuo3+LoZ7UJRm3fzWdxNO1NQ3
7DP5G2u/S6/CBoAfRELbehoP2GTYFzkZ1UX3dg3StMEyWeIO1aHigCrH7XPfh+zk
QqvRKJyOs3zBhdvWFxcTB+J6MFnsJNjHCj5T6OqJHBISvg3/G9cO3Rf8HIPyKi9d
Si84vsZd3fJZMkqyjPz3MtZ4+Y6/RAgnVE9nLv6dAHZYr6A8osyyoVI+EpI7ToIK
MtB/8uEV1y+f0gok3pwIuNJnzPiZHFSR9DvZdiFMLb+7A0qL5clm1L7smSePfZKH
D0XKU14+bscR2lgAgv/bcbl9l9YoMWW/JVkZ+uLgw+zmpn9HkJi9qGW4AF1OGDwU
Ov4e2OPloUuKiFZQI0WIfAdKPH+APAnCsULR3XT6PoHhZNmhZAHW20S/fUJJAqZ5
KnyuEyFrK7Q6pfslIy+UNalAUZhS7xHDSqiCPhQRTB8UW/un+oJlWMoyFs6+Roi0
y3ymC3Q11BaVrWUJaFtt7YlBbVXahoFm64Q1khuAw9Lj56ha9fQxmlGe2YBqN7n6
kWpw1Az4I97FXF3BoZbICf3a4yrN9++9mc7mkfjKdDR0c/8czehryNrK6je5uuME
uScqUQRWXxUjgytp3TY+hzyChgnDEP3OMuvtmPZ6z40tseZu0bb6sT3YMaMu6IrP
ktxsxA+CEJumITCR9pudobwaELMNSp6Cqwrf4qpRZYVaU59MQh+n5N4gmFkk6EBl
DyRbnOEUtnCk8gbbH3OZ8g1NLoEQrHR9+N+GmLjEBwMaKsKpmsR33WEBJ31NTB9t
JTrT20It5kufsBqpJEbsFvbOcYJ3mWLVgPuQ7U6ghjvLwf7glGiFhgvWQVQsg5PN
Wj6TBELC2fhf14WVSV/nEto0zGz6w50xfFf65rVITwuz4Tm5xLj6EocyqllBXOpC
0OK809mbgK/9vddFpENhzJNNXfkQJa/rK78JybeSnUgZizx53uAT330CncDIRQZN
JtC5GfLTkzq29Ae/jmhxZRVJW73Ec+a+5TK3LIRirhpyo5SQDr46B8e1cXMNSI9k
QHVysycIGIPLtRp49z0KjuADiwUQaZGTZrXRaiILzzH2wWuMUluO5BnvzQyEARX1
c7+ufnrI4WZIMKSXSJIVN+XE6yp6M6bRyJNz2qvocDDop3Ql+1KbpOI93raEa4bD
bI/dHhw7cnXgtM+zmmPkcBiKzKaL25iAuOht6Ot0o7zL+kMhtSgHGoFT77u52d08
CvgyTDV62eKc3fln09swuAPBYeVDF05vppDCQjeexMmjX8HC6rH6/Hgn8BPy87CF
NSWDfU5PxuohHCpHLVEWIo/XGyj7C0xLn777f0ojp6/semhoKIlPOPZDZLJyo3iQ
QBXCqK7fsujipClKpBPV2bcf4d1z0NO/Ilz1mFGs1XIosWiM7sEDWwpGrxPYNPx/
+JfCv1NCBojjNT39RdZ/Kp+y0KnvNvC641UUO2mVF4SMGIWy6/vRBtR/mlmf/Yxi
G4TjEb6UwlSTdXvyB5ji+FeuRWkRurHdhnac6BZ6bsaHWO7gTaEOvqpVIZyOz2YO
ecs3v5HRhzY6F/Qvmik1kCcD3pnbQpwNA+TsF3VAC5skswJodOeCF7mxO52rF6BK
Y2SeGkwgLOzW6bweE05BYbiOHvYLW6NU14tqkYsI5SUrjjqZZtD0HH4B4NZPKuKg
QRW362Acy2mx4L4zp2oE+TztndtQuPWDacjAYLbE+ove6y/LoQoLSxBXYw49FSh7
SP84a0XmGaHgvVIQ/6xfMFABu+3MXODw9IJVhMTU3Kj0Glz6mFs2guOAVfva6g6n
9MUuNDTHUtJAKhnWbd6RW/iNbUHe3+BXueEMqOVhm1FQdeoDdqh95JVCOeSpzly4
/lmsRp6X2w5AJSBP2HgEaxSMSaPIp1D48IR4/OVheArFZkgU1jq9Pt3ir3pp6Hxg
x2PIP4XrmxPI7XbSiWkgKa1+zugxmDhlU6CsV1hUGXqigtTbGsSMZ9Vu+wapngG3
ob+V2pzdeE91SpH7dKk04W82YuHFQdoU0lfL0IdVRrUdM0d6STYGz+hEcF5oYGDF
5szVKrq82KM0ZBmXu7kqKwcXg3mHcF6Edh1jcHqpps5FlLmpZa+6GUSmdhj/MdCd
Xe+/BN5rb3ohAokA1zSCXqsO9HccwjK9e0afeA+M6mCxImV+3CIk3CnSYE44LiTq
rfgo5HBQpzxuJRQAWmyzRqplP8f93XrPptD5jOmVHf0ns5WVIihMa32gHqBo31hE
JYvLc0ysadiYnWoDYF933Gq4yPLqmYTR1u+HRjcAxz0uB7e+uhhxpk5cvOEsCEbD
NTv9sBCYAsnN3Rng0owyyedydu7ABbxEeafZTF2tbODbmBVid5wkTT7APY64Cm7t
GZa17lKqrorAEpcPbPOaswyr6aHODflkrHn8cc4G02v8wlCk0NBHQ3Q09koaIsHz
L2Pohhs52rSv9cPfhHID5QK9W9Vk9cqJzya15KR4p9MXxTwyesniJnCP7MH+pumH
SOCzBgcRG9bfkwiywS0gD0vKuiL6/Rv8HvM2eOD1POQ/oZ7ynrG2NFScpXTRJice
9rrtbehBdiBMGx15uqeDuqXRBpHP0YYN8z0Hcb52R5pWFeTLZKVSId8zyfnXetm3
jtXk4s0OtWOkcjV863Piu+lj1icawiU3zPMHpzv8jrKe3lhY/Z50/7osEsG0iDql
HuuLznev/y6LvtrEuSsOGu1OdxhctCTg/mqhiF2DW7pco6bUndjSRBthZWyf1q0T
dyFQjwXCsdNPXcYcozD5NgpDCr+QW/iqAKFmrJnK1EpEB4kA4VNJrOOWccOLVi/Z
X3T3nZahgQpCS+rBU+hOiIMJXArT8f9i8lyJkdN28+vjbQ+m852iLP1zDTusY+oE
t6byeuw1ht1dtrqN0qcdK60zBFTfY3nsbAuFLTjYY9Ks0GSgeIQAd6T7P/lO/mzP
5zfhY+OnybssfVK7jDHWcjg1H8/l99F07B209+Hq5V34VrBSGPHcvUX95SCZSzOA
FhaEvn6bY9aXLRcx+phgvAlH000F00Y3m0p0t5msMej0qyDNSsaoOlaniCViE6gO
p2smWrXx1B5G8+SURKFaLHIGErlbkvPn9KI1rZoZ32zxckEbQVsWO6UOi1aOtobh
zna6EuNoYN3Jc4ABu6EAELegq0jml8waTIa+IjgKfTlZZ20moIs1b4Tf2c59sKIN
FQYb34VYmlacy6ikq2lBb+AVZYSLjFT48kA1ck7gFB1hysTitsW4AylDzuIJp8lw
IldSL5RSJNHFMYCgAimuaoYd6HfFC7W7kdwNL8+23oIFc2Apb5Qnp8baku4KunWj
mdN6FEufzTtbo11Jc/43EVCSXvkl5CLONA6ErvoIkA6rDacS+hhp1uufZGaOapxS
p6rwL62H5NV9w9h5kY882rbpsBVjQ2Nx2asycFGzyynOM6Zz5tKV+qsuz+65fBBR
stPlbYjc0Hun37fzbkjuYGfCNclE/t+TocHw/6Ol2LoZdJOTbXSJtVTogzawYHh6
7YI2TcCE4vPfqXcZamM4TNYyHdHACZcI/ofepu+SL79ZI8RciFvR0mBgojWpdmLt
rcdWy1qmz4a9zSMMgx+nxVABBPYUvWvYndLpmcpCsM2vosTzDRjFpA84D2/c+WVF
9CMKvUY9WrSkcJCZ1JdCRNPmLK2wHijJJFf+dr/wVThiTqxcbJuqHtkjqk1uN6oa
BQTl8rYi60JRawjZzaqX3aNGptdE0JUfGRAQoOPPAz57kRCxapDDbllQIGJmdLzJ
P83Gz/omyzdXtCdMPtGkpt9rCk6xlYT8PvQFPj6etcIpufVFn6zf6bkt4AS5iRvK
mrrMi8FcMsEktOSMqnO/dCbyFCmO91xfuqUADlqn+LJKpeJPMSG3U1BlKDmZUrYE
Px9AbN6JVzux8ePAdQDG2dBPz7d6EdxlpzOxdfn2onUagIKNbkH6nos+1KRTaNNb
H65sirbYpxFBpruvsYWHR4BgDtkl9/kK5vBwBqa0EfqJ3660I3Ak7uQ4Dd8Pf2vn
L1yze/RrQHHWhDgbIyeVax9A5bIrcxo66DwMbJam3DoOXWL7ww8R6A/1bZf0m3IV
vGLauGIiPwmtsUNWHB/zh87r401jaBUFgCgwJWcZFwM/D5gPiM1CR53yeNzMzhoP
30n/oi2yEwSyOlrJYitZhsFdOhkUQ0HhBucbxMFvo6zutDWMVjE9zMVKXamYYwru
FkmBlUjgy3i4rDUj06ApYMKpVFM6ZHgeru7AGZ/7fCuUE/+S1ifCjwCiQAIHcq7f
5rFF0JTKKgbt7PGYJX6lpankn80Bgxi0if5Hzax/jJasnQDW7XNdmdNXVHIHu6V6
lkRFxyhYBNisgRCKa4i3pXEBUVsl0wGuZJhKhw98kY7X7giUgw0PN7ch/yad4g2x
2BDJj1062pcfeqjdvvyhtDFuBC8Jyh+XECPJm4CA5Nrc3OB9IWh1lf4nYuL0pB21
9GQ+NBoLW9m8FdxFzZn0qRnlWGramRG8otlbaYHJy8zJIZYv0JgOXXZIAyfsg56l
L/9yvsbiSOMBKW4ocz41G1QicioKMqzb03cmldjCBgPX6MYH3L2GBu5iF0u9UobJ
DI9jE1VcRL9K39SKHQdBQRqJv1L85zWAr2xn0m2+ORLZVicfiZZFCddA49Rn/lto
H8u0sDTOFfCv/FKWBX6FXZg0XHxXL4qQAItNyAlaQ1nVim5vu52MDPufE6uyP8eN
AwSSXcbt4t2vkL3Hh6iVeG5Ri6Qivr58nJ6U+ZJBoiMMgtUCH+tgCcwp/FV14kci
tjYcIFJxd3YvXJFKeorgr+TsuHtRQBy4YdPcyCekUZM7eQIN9NJA4kM+XDCTrB8d
TUsOYTu5PHFlmR65aA5VsKRwr0ZJrQAvofF8bWcYFfccgCek6q3tPEYCPoVuOEwf
eY7dA+fA96d6QA01FczFXfTDBuoRxKvrrcaNVWhVCH2CJlPJ/cHvkc4JTpDlobXJ
PYA8zvGd2/LS8uB7F36vHJhlj8D0KhIxUEeaFp/jt2CLZn4YTtrr6t9u4hXb3HP/
st3PyyEzAs/p0UoSbb5DH1WhCjeMt90Lv7LWTSiM3VBo5Tr4fLo0TGdX3y/aK2L2
vpAYrTnKcYAFZ0Z9ch6kXS8IpnkDxcK3O3s6Gi5LUc2UedQrKlVUHPz/oleK0Ogz
iL9mqhh0Q2pjVmUh9qZqXW8AdWJ7jNCmI8V5Q4TP3ieLUjkfTgIsbiHZuUpS10on
eIxBngW7mvWCzCdXbOk7l2M+5HjViJARhYIcj8pCxJ4SO7Bl6rP8raiG6R7NG68i
jTXJnTuaMLIwo45zHjt/TD0A+aGQmUHUh6eV0SCYad+Ru0Uk51qudvg1kU+xeUfY
Rhmm70doFTzfa9jO/ZpSV7qlsGWe38NKxKErCpjggBUnA/aWvrGPgI3bBoKYsdrG
TkDODnmtPPreg9LcGCkFNvbngaveZgNmCBhqOs+eZx+GLlWJYmN4zhh5mNSRaZL4
wC+RI6GVtL/81MhVPjKzx51hCeF1lzfB1I5uWLhQaDeKC0R7lhM8H/fiBa8PX83z
EJGQ7sSZRW2Ia4m5SKnotKNFL8SCCs72eyaL2Sqv7RmzVkoRYO3/PbCrFewfA4wn
Hkwp5gCjYOr/ycJ/Zv91ImnYoTACMR3lSJlHsS1H8YI0jshoIEXABPTSUYSKzTb/
hKF/QMykPolNFencrgXaTl5U/95S/13/7WQLFZt3G3gzSuQj8FopgGocNBLB+ggW
dfkG55tBCiTHtOT5dLzcOIgntYTpJRUBVRsewTz5DRm19v6Iv38e5TjCfmUcpjRH
AqUhkl3fENkW16jR1EVhW2Yjp6AMkPrT2mI8nzYTuM6i6CW/K8whkccH1mlURebe
0/U5iseJs80hOz5NsuU8Amv1/FFkjEa2SpkxWcE8OfU4shYWXmR1oBR/CYZ9H5KQ
Za86VcEZ+lHED3t8qVOSrligyu+B/uA+BdSa3v2yRy1YSAz48g8Q75FMjxRVCnEU
235CZD4QtXvXR7AikrBEWFeh9MKnHNuh/KQqAz1UhfmToz95ppLt4bNGBOWMhj4Z
b1plltL4CTm6vb3L01IKjj8RlAAHJ7xXqVO+W5rwHE2s5+FDmNN4pSOx572U3MTy
pdWxCMpL70o6Dvmy/np7hn6HF6esh0i+II3UT1wfsmyhF6EPuCvn8hXbgoCvg4WP
FRU5btFznXcQ3+D6Wa0sNVk+CBhmoxDaXUoYOjVN6mKFPezzekxY1h8gCXA4A1r1
fAwA3Bg3vmVL4w54P5ihP4Ypxf93a5/QFOqXICpRs7bNfMTB8QZUDiickvVez8Va
jjzKZ686tsip3I6cQuXYgQZ8KbsaWp1A2Z3b742uvsx/yuenrlP2hH+VtP9PY16g
VeNJou/JG4KPfEGX4vtF6e/aQnOpf0dH/xiLPVfI2GoTFqZ0wqo8anKEw7TG2kmj
0GHzl4cHfugp62as+klxYtP8OBMtghmkijKbf6sB09tudWor03ySHjETZ+J1iwPc
Mw9tTwv+2tPNE/nKq8v+9WkxqQ+C70xghZPIjXM7Kkgl1BoUzkgHRhoczPKAsbxd
s72ACdTDacPaQwcqr7p3djpt11KRqytUuPLDmkHctnIya4EUyPm00Sa+xyT3oScj
ryO7dpRG0SC+EbZ/O/kYTLcN/uwlFTaPCItuNSdd6YhLd7XuI86gB3yZjc/UAhDI
wwRSeISBEA5srVH5A2fuWcHwjo/9s+ffc2SRmxMvzbz0PnnzrXY9XTo7gT6KcJDT
aaR1mpX5AIh7Et/Gu3sH1Ucsa8bj4urF6W14lVacfiSVPLh8gPYEJfmXp6pxuyLC
LnQgcpjmtMAltZ5MTkcW4pSfeNP3ca+pcEzJP8XZU3+6L09VlalOjoV8KmVR4//u
WSowJTtBdHZ0cajx0kIkCd86HZfnPZHP0HH0Vyt/9P17Yx7pjZYNfBFX2gLIPmTX
D0W0+65prURNqO2fp1awPQpv2gEasRMVlxt6YO1bJKfFR/56QaiShk9u531o1KvW
pt7BCm3gDO9jOftVo0rTQZKRvqaF/b4SiCCRdpk6vzfYCljKDCmP6D0I6LXPSmOs
L7SE97cmDCs1deohWB1WeDprRv/w7YbbyEYjtp3VHyR0tulGWPEpD99vQNJRDt2/
4dUL8EQv5Cm4WfOPlSNrnBaL5sBQjp0sTw2tJpFMXklk3FYP7axFZ+PU5drUExZ2
Y8vhxOFWmsXyRLASCOMV43YyofvpOb8yQ50vTvBcLz+OA2X2fZqMgUHYamqQFEos
ZRBynlOTeZJ+MhpubOFqUL2PCs1Qi3sWLfwIV9KSNyMVW877iwn+uQUbWWMpHi//
lG908WZu0QTnVU5dCw2B9jiynX+N6WHog8oNFRYAwWwEgQOmvZr8EhWUsy/AAVhg
pDEecYWPnwNjxKJQuMk1ZY2SE2Swxox3KASlbfrEizWQ1T5iCdGt1L3Uw3O1q4x9
RFPH3cipvsfh4F1ahouQMFfqfJgOx55AnS6yGbZYIvZ5O6Nu/zugbMjIAINxI8L+
wqzqKNp1LET2pMJ9pRDX84LLAyLtS4QgRPYeOzt5PDzFC9w6RuWX7XTR/vjom/OB
80wYbycQwQNTGPic1yMvTuBQiVKmD9088fbg+ndgPrXdCAr9EQlZjuc6Mxfki1Ix
JnRyIBWK/Jex+0ri0TnWc3UlHLwCM+ingvVZY/PvBh6NituBlgbTHslCg3yF0WOh
QS3TaOjFG3E3ulVfVp10HqGHC3MBkwZhjul5pwN2lk6+UWzTQX1Wy1mWU/bol6Ie
7ov9Qwi0BvfFUKR4JwCKMoiLm8OJztVF4DR4X0ZnMsobeOVdDAjSR7oM1w8buwfn
1LvNq5CXKL8wX7xwqk6LmbwDEjMjkb4pLbyLQX0X7koNJTd8vcRKS7R/8Zs3gfT3
Y5E/QozBlHAEm+OOBiaRxNSGGDv2CmLKinYzYGdesW2UdkmvMmW0/yitx17SEe6u
4Is4wg+hCgGfTtDLQTZV2PGW8jtH4rs0tkQD/gopRz1D68bFNHt8JSmzUxC6XWJ9
um7oGZerOn0QGZXHiikWF8tf8WHfdQAMHYQagKsDMJiabv4o2Dp4kbm8TtR74dxQ
B4KNYLTEOyQ4e2cgX21eVAWcGaleQcajsNOmbsaG4bwKFkY3mPqfJjFo3HhYhRAx
Qm6LH6G7cqSce8eE9qk+UC/SlKaKIaJOOc3A0Gx2m767GVYAw530h5Q51vW9AuxB
OXTjFr/xcL8BW22E2jIyXEwxdYrb9PMPGS51H0cyjayvb0uELiDkwJDFZo3wy9cu
TszUmYDQEhhTGKPGBmaHovVD+4QnKy+WDZFWRZb8Hme5ThwmBhtRawLb+R9T3+3p
qYO21X67cJFamgrlAtpXLmOyMSqFEC6Nf+25N69YGGah1VqqjHn2EEnz/qmg1LMQ
uRog2ljgkI8C3ioj6wiQLmpXma1Ynq3NBpgshnw9SyRpxcbKWTPeggfsIq9fja3a
LEm2cfI96KkTx0yukOMBgdyqvHXeLYUP6Ui9VfQP78+sWt6tXMembJpG+KMboeSr
Nsiy1abtMZOSdoC0KqMArczxAiLzZdELDZvRfGP1gDdh8fSjjq6yEIuhr9FCzANY
9rwkoOSsfqUkzuooE8wNJY822RNTEaTtsWmGzvHdzYkC3Kf8HGW8sWLJPspuRuKd
Gtp3r4F5/egB6g3gRqfbPhAOaMSU2MRlgNnVhJMK5fXMlFmE3vJUeZHvR03c5v7H
FCqGkyG4v764lzsMqRw7+4yZgwU3aHCWdzdjm/y8F2C0EEcNtvkf087g0I4LwtCG
9NMNzauVzA4/sLTQGAqO9gCuI15pB0FRdh41o9Gna8f37OjznzXxPSVPPjjYvRw2
NP5AsyITBYBOS7YrC+nM22CHYkysI0wKodNyakJpcrwM2oSwDj7Vj7T0rswI1BaU
L3sSU7u9M95mpYilQEZc0U1ToJ0A/kWItaGzrD9uXnsPynDDHev42lGDPDGetQrq
19XWT+5jwXWBNvZs8N4zX5hXrdddekuxzIMJsOW5LqOCyq6iZiN/M2saU2QzpF58
OGe+RNt2Ju6Z9oyqlwrXnk+SP/xq80XIQE2AlbYr3htFStEIENSWgGotLW5jdXwh
XzBvoq77Kw7AGi3sdZJlzbUax7z2CKkfLDARr1t/5P6rnPs7KtVVxlL9eNqlz4mq
DHTvljXFTKaiqil+D72b5PNNM7eND5KfUBcr6rlreSPAAMG7aXG8IGwX+QKvKJwK
Ao6Lu5iOjmt70WFCrn3dbkJYBZ/VE8LI1pP3qG/9GrzR7jJT29pzjl7Q/bQWn9rx
F/S81od+dcJhqDUbmj1De0gd441w/ADM0yjgRw2E62pn+73wjSgUsjKnxbjeiyJE
LQoSWGt4ZHh8d0Wx8zljavrHF3xdo37tvo2HRRiDBE1Vm+J9SYUuPrTypYJ5doIG
MYH33B4GWBvcduzhl9uVLiYhsKGhPttRPFFx5qB3Xqk/RGwcikin1M4llJflP8uT
9NYlAzxPWlaSHhSjXVMfi+S056U7Ed9fVJenk0mdjCIE/9okHtbkPHsVra+yh6oL
g+331m64aAwG+bw9+QM5T5mf3BaCRdjn8AIjIi20Z6kZkxtFEbBQV+jjNXiy3Xot
zLf+QpAQqgoFx3j233vFdEfY10fRCoARon3dlxwZJqdsEAaih7VaTqnU4MA0dC/f
1zBsdnjixp0zFBw32eQnBAVLmdS6HldMkn2dC6Mb0sgv3XTUKg/CvcRTyisVeK4Z
pRAoXTfw0Zj7tDIX2SR+wbkCLrwykL07rFhrDOoXljubyTruWE886tqsRQ5k+v7p
SYDVfEDYrurhLV21eYDO3WkIbNXLnvHUhG2bTIPEg5o8sv0wXKryg70KeSroqaU4
TgA66cFRZDSc6Pm+kfwUCYwIrwkT92za70NvRHCzUtcyyQ9yOFsyKdcCGsCePkas
U7mA8HfXF4MVrMe60bRjKu3wL9+k79NzPfhzdPepuF7IOCo7dVQN+UwyJ2ib0WdS
nq+shsGyM1z/LNtGC5HuWK66zeK9FKcXRLBSBHYbHyUHyrfRF/8s64gQ0w60/PN1
dzJe2Jfr5q9xR2xP5s17qgsxmzA7B6J3iH0Er2EfS5sNbGfQ1d5qqFt/dc8+QTSV
fRW97Gg0KjBK1sPFjwFHv31ZhNNWpT+FecKWpSLBCrRlfiDIvRvoPrj1XSBR/yBo
tW7se7wWOG1vhh5ZuM/1TXF1axHgU6CM8h7OHvQDfiyf2bO7gEeY8wWF7gkLJdzt
gFfRoa8zH+nZa4v4xpCuYvl9I5hpaeYUMVky6YX3i5AMzHQcfLFdnclSl25REgqM
7So2VDNzILgVlTvcivkmVC2Zcn+y6ImoYrJG6DTswGfX0jum7cPvl33rVN0KenPi
ozIFbQ4Vn9lQ1AiGBLlJqWjwZGZZEh0/7ThV5qrnkFQ9lFz+y2SDgwbtkIlRk1IU
xhKcEeKsU+wo6yv6ENyqjn82OJv3n8qJ9JTb7o5sAW7YOLTfwDT0wJN2UBTkTg/W
d+Vi02N+Eqj3CTzoVcqNzykoi8cKl31WU1KwUvtjG8GHhluYevCmnu7yH8aBwuBr
m9hZWwNZDGoBe21fVmOfWBPFev2QmRiG6wt7S2K/xdTvZzht/gjx5EEkTNPmN6cr
urEX5nfvtReuzCIHblsosXre0N3aAby+pfDMVcnJ1Xor7HJgJvsm0RZ7vR5qBckn
9kRHL50yoYQICaFusX0OSguHwT5fo47lNVe9kY25i8LgiCt8Mtq94h0LmefFKI4r
A+WluTbXKAzk/6M/fZ78Xhu3+XTwvDLXc+8fq/8yIimNlPpAALG8+FWISGopExB5
ZTG9AKW7Lar5CUwtrP2XhtJxIpMjvaNhcTXJFKYrj7DfF74YtdfROh/sOT9iBRgm
SHwnpOl5id/Ge9PrkMeyPR2RMKABpcFDdVpwLIjncuUYxRZykn5OLd1qJUjzj3oO
TB2sElJkG/KxA1Hj12D996d6ZNAbFU516Xlin1e3LCGngDL/xQpIAfXEdXy8GCef
CGhfK7g/g0u2de0v3sEtyfq2/cM5rM+oMMWF9T5kHnU79MvVK6oM9FzwxsBvo4QL
s7NrRVpQ1vMK24Joq+hUM4xknYSqKarH3AE1ZEOgRcDBvXTXhFbZNRaGxsax4i45
i+i6pXWcRTZ415MQT4rf1O55DNpcdVPonD+NIzF2VHy6tjwCbsY/dZxvyj23hNgg
AHz8iF0j6T4wP66G0vrbH+p+IizpMIjsdi9MZ4y5W3SaMSeAVv+J7Xt+Zr1qg1r6
ilC2GuHi2UNG10NczBkkSCyBnhLo+StqNZpK7JPodjDsf9CziiqDtUSUH5GP4dHC
kibnfVUsIthZM7V5ogpRGwFniuWC+gGZYkC5k+z7lw6ciBotrWc6ANe3hPdSw7Hh
ksorQ3oyiLQSJn0C/UCIa25ewtY5HMFqA2C6MdpWdiYuJP5/vx+RmYxoVwUt2iad
8zEZbazqV/aFfxYAkquGtOuy6Vd6sfpSRyiFdhb0MDX2Z4G4VadkkJQxc3gwDJe1
VEadp66zMqzE8jnN0C04qYx3rWlEnHL9NA3weksZyb2pm8NFCwVkCfYwuPXWAiRv
ydkRWoEkYNtZWyWAswO2DFREeMzmUFFxDGZo5/HPCCf7R+Str0nhppKKyyS/2Nfj
dedpq7rk+DIJ3rfjqNDjN12iguerzVvaA6aTvq91YRPxRZHPO6nlxAXObUVQqHGa
akjGZc40he8xq0SnjFGK9DTsBDc9EJFDpyof0WhToe6XvSRULiEr15z+m8i/+Afl
cu0uC16zzw4O9YGnFx/tHtdTVrEilFDJLEV+zda02HssIidL+i5+S0sdWyhlfQ2i
PqyqaJXUkfjm1gKlaJHXBHiZih7O3rJ6sXZ+XIum9PtzrTfvixnC6+OgToG3KGaC
9VDv/eZxXOJCeMCWkdHrJX6Pf6i0+6A+utl7Qf3U1qe6MsBkEWNPlrtV5sV6urKy
BnMUTczSMUDNzN+s8sOySbfjYdxRnvs9tHww1J3tdoZDRH75/Db60jjs/87/zjxw
iant1fK3JZV11YYKmIF/94FhXrzzajsm6aLFh5rDgGiIJGkdl4MpRMXwz9qdHvol
1MAGJZRjn3YIighEsFvX05I88CnfbSO0G0IyeJemrmbXDnIxA161hsbWcudLoXeJ
Y15yOoJZUMCskejmXrc2lhdULaOszx1kJ0qlv+6IptZxliiSI1K5vfZGEOJU0+eF
ballrSqQEG3eMHphan7uCGowdMhGQKHgobJBHqkJxwgcLAK2LO98YaBOqGTln0t7
bMR/u2qfKmihUajRb/pn9c+LFCqirEn86zc3LyQy451A3C2Gk/pQSYEsV7tAzAt0
uvAsi/W0aIVPq1fNV0qsIzxGxDmsP/V/7gvcVkFgAFxRzDnEi+MdUXWu0d3lEnzk
kTfZa3HjPbmlnfB5sIafW/N7MDTMXPbeFPAJEHFl8M7N9XALc8vSWwz9MDRBbafa
yGM+OT7gQ+pSsRyZUnMoLXCv/RFjTCcifLtoT9TZTQeZGU1tNT4URP0bQ/0rj6CB
0R5tBR1uVbtOojCdnwMd0ntrFtJFkTjKO0OER/MFj+uFyDEgtGEuAetd9wg2hSXZ
mYSJO4UZkUc0syV2iZVaqxKmzU0zam5adXsMML9mSldzDWtYv2xqvb30+rrBM5xb
5jNfmfwmbsIoUObNdhVLINt5kW3rk3eKppm7UF+BiVkUZDRYJxtTnH+S/HhoP337
dvWHNNPF4VDjVOeW5pMjGJatDV1+zWJEs/P1KaF4gP8N007FzZY/M42sV6C+c/QQ
mKEa1Tm6PcGRXG0j99HDLiMz9H3ISEYDCowgLjHeM5NunDplIYH4TafEdNcecOXp
RCq3xZMIwznNngun+g0mbN+Evl943YppeknH+8q4oHhka35wbGkRTCf8Chbc5ihk
5DofSr6DZ5T/M0xD0vJCFGt7P9zNdpJJmWzF6ZxmPQrupLAHHbSYyr3nG18VeMKF
tjAaZ0z5DnzTAsv3Rt3tCnb282mpH/oFni2/68yzo8si0AJKND9rWkfKBZ/JuPWd
bGuEmF4cAzN9AwOp/FgD1iekJDrLrgzo0V4OuVcXY/XQYyqbJrnmlBEebz2qOc3Z
LifRNsBNplCspVwTnRqo4zrcLPfyACforv1WC/VzVKawW+yFupaMeH/i8tTs0sRC
AQfIIGIxSFBiBNRVK2XuF8kOIoSc92wSxXUpfTFQi63Gt9Ny07Q6Rd+hDzJafjyz
BfwuymTnuiDPOdM3In9j1o0wePMAvpYR/x5hBfSc2isejUpZ6BSm4y46Vov8dFbG
1asG4XDTNzMTCvWVQxMEjb87WVBkkMo3sjAQoDnDpSBPXxF2eLlLMcQvFWL0p/bH
cbaIMj7jKX2VmaI/p1Aae+KUSm+CwV9nGdUUdnmQ7/GoFwgKrj0ZXPt9uiO2EKjc
NClFL6o0duM51HzAMHLvRf47hvRU88lM76ktSFvxgsAVQKc/bQBLqMrTKcb/PhZT
DMsKSPN2UkEecxkhJvrDdUSazC8wiij32Vjnb0USzK1TfhFLsblEDo6eCrz8CcjE
9+f3rKw0jhsER+nVbFb2HbrRpLPiBqpJObjZmbPzif0S3sM0n1eh2aQYdyFNqz0o
WD+s3YNyHcSBV6yvbg2lNAF1eEcXT26BVHJOVbQoVrCbRpyfqY8fh/4fPgc049yd
BUy1EaoCCNRqLBghOsI0r+BgIz+vy3vvIIoCve6XnG32CmkaRXMJPSKUb9KOc/k2
fkwqgOA+sKBradbseRlKVwf6ssgIoaaN3PFDtMeFqF6nZNnW1eog2ntWhk2EizoW
SkHfgFG0jDDDlx8m9kl1a/BhuR8D0rLNdU9Qgn7+dRGlpq9rPuaCZi6USF/QhJFl
XuKqMNmlzjOGPrvaAvm5nLKbbXZr9ReuDH3YZtjdHkujCQ9JNLrIsIa2jEwa0cBY
z7B3gAA/jqXGzeNPxDNaGXaFERVLhNUKuXCKk5eeRuxB/Z98wlze1V2Exas3hlyi
BzTAlkhNv5d0svle6hS5yJn3OnTxFxKJHaU9756g8HwJuje1ldxNqI+c9g/Xvv+2
Hfmp0WAcgY2gX1bHKrXysk8KgRItgQWQKQbg3bG6zDS21tnoCxDzDEB0qQEpha//
fmqMe2aOKDVgTbUlgwZl1vncfrDbkAKMMYgMlwY4QCQL/J6/JU9/Zosqlic9KpS6
IrnZ8uBFs6OECSwbldOwrCu7w3tRmyhl9jW5HEnZr2dtzbh/qcp3MPIDEO6kjx1C
CqeGCGIWAZB4gXS3ex8VNHcjUwUmf14kzepP4ZZ2esoGbqyIyM4q6cfhTRVjLFQw
FPk13rZKlp1KR4gU1sfTHJ+Ac5mPl/vfdQH4rpVB8TBuoqRODSHrz8jeBU0ZTqtr
IM9Pv8Op+m3UCeKPC7DX8sPRh6/5tSNHRDxkejOeEWiLRm3lpdO+ydlbi7qvrJcW
kbCrKgqYGCRnxPwyZ5yrvIvORJZOXF2byZsHnHiVtZsqfbAgSiAcl7dB50kf+sMF
BskZYcpi1Fbk+asA6cKpHdFBgNycrRLCPBaRuZnnHausgh6iLgDS3LbWYmH2fedR
tvMpT2j9op1zEavV3h+1tU/uwtycXSNOCtoMDCUmEl5oBYDriTTaxEeyfGW1OOk+
78vH0BeL1Ggtouv8x4bSqxo442GFfK+AeJWALxq91u1hIpUo5s1qjiKcIBieuxfL
P6Fs3j4LUn4t7PEy6wlbGt+tSIjmg1t6cJGIei/STG55xTsd+1sh7DBpSiD5RX6S
T40KCuF+V4NPbwyp6osWEyppFTN2HT14WpYDNitZVNhvWztYTYe5PLJajvcbGfGz
WMa2xMMIpS4RKRBRzm0CO2PUYsdrJYznmu+V24IrbDgJSngF9/HmH60eivwLpQhE
GhEUo5XCnd8l8N75Va+BSAXR4RRKmdM21mYABgiJDjp+5LcJnf5jD6fztVHRpp3x
p2C6LO3zq+M3E6vHsje9V0xHsBLPpIBAqNgXRHLnP1Ka9r7JhWI0loe4EoXP8kA0
T4rxnntWhpMfBwm5WAJCEXiKchqwCXe0/7aV7Z/QLxsPy+L8KCVaDEhPehimXwaJ
3+6Vqo4r0OEKxFzEONF4mf/Z/6yDKSoeEIMaPrvsF84CAyNnV7lRJgPq/AW2lxfP
9oRhyAdFBo/u1w+dZdwet5KeHdwUrUbrOsghGfhGkMdA1P1CnYkFmtRlNAipMLnN
EENT4X4n/saH6srWSlReMbJF1gZrk5bOXaRxlTQAGZi5tEGPFhfwxcERzsCET95Z
s67aK4DSFWUVEXlSveObDiXA1TE+3Gg1/3v+4WysBZdiNkCNjQ37/KWFtG/cUiGn
blVLMFouZyLdWami9xYefVVcijHzQ86Ax5xA6iVJYtwzneQ6rtIFIGxxbo/IEmjf
0Yj7dFFusdhGj7PTvZZkvlMJXgzfKCOCVMgzqWeSf0RraeTXfQeMHkC94ZHvH+es
x+9Um0W9omoUyNc7XvJMeVuZgmmWOiY2yQF94Co2Vdy16mhnIJXrGN1pWneeTXkK
v59t1Dbut6bWxJtxvDl4dfmiucGhtL5YF/cry/nctv75f/mWRzrQuJSqpotVfNmV
g+8kI1Gydh2J8acdlwWWAGw50EAaopwu+pQZLNQxlUQ03jZplHYWJnPG506SE0JH
j0XJ+R9bTmpQ43NAQixMjzd9g+k52zYG5HqBbdut0EUzToEVIYk6Xwp7eVIbnXZU
AQeZfXu3V41r/DzlqcTJ7grPBlTVVGsQYf58wlSeoxQNdqmMEvU+ejlJbgDq4Vhc
P0bNxQ2j0T1QJCspaBYVhmtPwTXsi7NT209k0TLMwCLN8MxLDkH2oA4/qCiC352l
9pca2GV2r/bPOvoFcoixFWybGc/92iy6IpKyeA4NaVgLg7BnuSL4+saI+Ut0A60H
Do8WTbtBNy9s7VKd8v4M5E79JLJ7KQA4WIZ/a7Ai8KV3A3OIr4h+TRVjqp/1k427
36f5UU3ZNPvTk0e9znkpZNqFD5ntvHVpaC7zgxIXwK1mA+uWBVyTV7qzwDn8JE5C
+jsj5/bRcWOPnQpygYSQcXRaBuR+rvJEhC21Af0qobE4ZuJv+l32AANi1UCBFfhN
iXdpa4jTksiWO23w9iAPYL24vqGypwCWhQApJ+p2JvjAd4rSfQLhf/oYc7u2OGqt
Nu8U8pQsnquh9WLrtlyR9hIStoDr1mAe0kEJDyC4vmdo8Xt4M208nP3+2g8dgbAq
wJREz8ZdCbe8nYCepupe5zOnyIqEsMXRY/MkYCQhQjguHLLhthuj2p83FpLb0sEe
xA5DR1EFp/ZfUplINcIId7HSIhyel1e6WrwdDvrDPSTtnn9sHr6YXSkNoMzD0awY
KeSSfKdcVZoKFaAwnB8It4VwUwLTFEy0VyGCz96wnitQrX5xEKWULITI+OTuhByt
64nRTgFx3kduhBYrIMKdrBEqZiqlsbwgXmNt4fiHKxhkXMQgVgkfgUZ6gT/6js6m
7Yc8wWjV5DeOmOSZBZc/9soP7OSNJyUgi3cqbkcyCmmz6RgBE8KUpCdAQfcnLbP6
TBrVDV5w7qEFkHlzyneNIW1DL1FQjcecwmwXN73w8Iq0s7qR7iX2AcrGiN0Vb4DG
ML798BLxBDioLpbSB0DXNe35GsAJlLXj4od2iPdeElwybFCTc1HcBy7H26TiNTW6
QbizbQVUQCwG4tonBqkqr9CcOaJsLiUdco+ieBT6kVo9tufb3FHI28eQipjtpw0a
n2ujqOLvnUSkCEcV+fCoY6YsD0iHVVXFMzh94fg3k/O6Q42Pk1caVp7ktJn/zBtQ
WgGctmr6aY0cOESlP12+BIf+z8sVK6wccuvVNepCuxXmFjbj6spsCoON0Oy2411w
WEvzlkJFGwP2ScGSbsJ5k+CMiuA1vLiDdtwXKP3cFIsBAtoXFn2REl9/ni2PaCeQ
bEG2PHWz88Jr2l4xFCrJc3h3d0d1JztnsygMa7S8WyPLVPMfbY02A3WBIMDYZjCk
Pxa8FudvVSkzqQsycG97kIjIYtdOkMbuKTm2WN6tzglOC/YfRSwdZwvgL2/gseC1
5UviNINJNts4AH4eeeJsXbi1eAcDL6GIbQ31X1Rh9F0x8hJkgHnZbmWddr6w28TN
loD1sddVvDaSM3eW5zPeR2W93eS6Qn8dbyjbSKeewf37I1jAuavX5GXPgbPtXB7r
ARH1FKBDeSKNXLz8VItShSSpI4P1qafT9i07RsgTA3Zqs7VIk6NBGHJM/+d7plVV
j7Tzx75pAQWIz+jxQWmozyqteWIIGuWoSnLMzoZswwBA/wP8+jGKC+ZjMi7EgOXt
X2kmA7aK0B2iQ8x/nZn7SYzs3aA0rUZDnqsAdOq542psTBUK+6P6ulyQ+0yLSuh2
RcJBlHNfu1rGtV8IwlB3E3WSovhkYS8iwU69p4NV5WDMcNnaQieXq67REA+Y676s
z8GxYLBus7T3maxDcOXLURst3v2xhYa0OS4jO0lDtTq6G1f0KjklytyYYPzRMyXf
i2JU+dEBrCxr3FCUIhLiHvarKeR1XIFznEMMWL3Kq/HRyv+7sNyo4YDqQ1WfAsXD
AaMRsoXRpjqIy2fATBSPsPogFaWwvFInCWjYVj+DEE42Rd/ejzwwwZ14Wbe7DBef
clWWWiGZdhFE2UW+Va8b9h3Z2ind9JaPnko+y6dE/VcFjacHIrZxV3LcoTi2kTKE
qaa1vNkgfUqTUWvs45Ky3di7QDkKGeEzPC4lDtfivcA8Hhr6hGirm8p55R2YVn98
hGDATybSeb7ndVk92lR5WSwIuyu3plYqgOFznF6GQgAbP3HzfO/VXmKGI4sCTmE0
RidJY8yMJWXx0HdMb5Vi8bCTzUHj6JVPJJS69csTGiZWqWuoXiI6FcW6AZlLSmA7
WHHyjxFGAEJnDNv4qm8C+0qbTUaRD9jTbj5/pJ9l+gNEZNL8V/sZO8y+B5nQpcS1
VlF0OCVwdfnnbFusDMTby+1mgJlbcHmNuRvK+3a3C4GTpUALSxjSwQH/W8L/hFso
4JWCkZKrbhmVU9pBonBEsykUiFaK6wlXFzywt5CtdXWGzGxsrM50b4fhXOTrIJuE
MsAzIxy/PffO9x8jbw8fW3KUiW52jswyvMaOfAKGDZBEWV3Sb6SSoq6z57fqzEfl
vMwlhf+E3yfWOhHZQwu0J+LktY4b9WGea6ABbYQdUF4+DRhJUqSxmxkzPG+kq9++
eKAbUGg6+jbkOt3WOgTQg9b/FYBG5zY5Vbagl7ISZTD2dmBAoTFEf4+JS4x6+VNZ
LeoWwQTl9Tu6F3b7yVeuzUzbGjI6gSVk9EEQ2tMKl287Nt9JU2ifumxQTkdzIU2V
tZZM9g0llbH3u1VIR6mm8s+mKNncpfnEkvz09UH7uQtDlcZN6STmBsr7JZiD2i9C
juvR5VyuLh41jEqaNudIr2K10apa6lvANDxjRDFXwS7o0dbMlWKrH4by3XaS/UFR
sYTzF65N9r5yTcWgmQ+CfFugUNEdFTU16EsTnNv9Z2Z+3JhkVZNWoEFhU2PBg+6P
DDGRJtjGLEsSpfxsnvMhp5NhLnbPc9pQsHpi0kR07sLRS0bo+eFNONZaU+dIEmP5
/CmhsRdFiZbT7uEMTk2yzHkqwFEB+uIU0uBk7nrNuA+YGRIGfKy7JTD63yX7PA5j
C6CJrHU/esyICOsXpKVdSMhNJF/3dUXVkWsxsqsKHHGAyokO8Q9gjM8yLQ0ZP6Wd
tUrM5+nviLgrahUZ+nHUcIyJBmUzaKzbg/X9nw7U6ztjtPQtKACXAE0lbWASit1O
SaySSV60BnSBxB+3dYrYBsSaog2k80XfKsSsH1iEDa4JlnDdSEJTF3X6vEZrr5Kp
QAXt6pv4XpMZmeXZEHj+9W+RJC/usjtpUcO44Qqv575zhyAgcVNJcOkO3Hs3JhXj
kHhieDgkju82Oqv2QrleREmDhPjIeM3HaIpMCbN1dY2Tzt4UklsyGbmw4jDmrbA5
e99vebKZw03OsZOzb7Jymz/m4sLvkTT0jxrfYZEZLGv/zemF8EEeZgutsfztFVKc
roptxLBZo6xRB1mlkYJB2uJ5AUEjQi0Re84e2YMPHV6T87FTZsnphCzsPgdbEUxq
m29slz0+zR9CQ8lPOqnI9FFgZh8wCnz1z3iS2TAGzWLJphAUcqfvjAMJjaotM9/9
+d1nHCkKHQeVDSXOTET+FhL66/DAZ5Mi9WPfs9alWVQYHtteOxzh67HOH45u/0dy
cfK9RmBsASIXg27AqB2onJS/yvGtEf28seyqI6aAH4VE7DBd2muN+e2QS9SkRrtL
6JNkCElKRuXkYJOe0t0xtk9JPja3KIrWJQfjn0qYUo0UTD+ntwe3Uepjff09asTl
XMn7v/kjF8uRtSg4g20gvCDrOTCO24bcg5HHJbi117zopm73X/dceg6LtI8JHMpr
fR8iUsdJ6oJp4bsLO6fy37qRcs/Ug3aWTBinkR6PeRElYPTbm5XbDd/A9Q5lsjuq
OdHsNbiAnhabkyr9RmYd1a2zOhCalR9CK/OdFUv24km0EWPG5if+olxeyNrvvz86
j8kL6SuVFy0uDlIPXpQvPk4oMaRPbr0XXZXw6LW77h92eiihQmJWdVU7kkXFA3Tg
O2xd9VP6Ec7A3WDDw1Vl6DzONVLh7CrMs5GCk+SzY40QS7Yf3/7uHnnMqKxL/BuV
E+YFN0V8Q3tSWV1/FW0NL+fBiquURVav5Ootsa9fG/+X6cUW5dcuOiW6qLx1gc5e
uVBhYH/sINggmckohcz7wwuNcbmE/f1NHDxzy8kQp3M0iBVxl8rpNXHNIogItP35
YrEAmNMdT/5knXlrH873u2tnJbHEgjqOZCJUq3y/cYn468J8MSLIPqGjAsjZJvne
XAjyIYSVyY2I/7jkRAeVgRFiyiGZoOxCHVqks+xbsRemYAiXs0DV6ISU2mTQsfjQ
M0ApBup5csjDHNJL0Hd0Eu8HA3vM2kBErEWA1VCtbgwFA+KP1eznfxeUDANE4FsM
74eVmgiqeSY4YrWIMHIK7TPXyzHd++liccoDfkoUDgNho/czwa2K9/doKdQGXBOx
TdO4AOxDMw50EIghxHmp2SbZlW+KZMsxFD5zQhXl1W1a7crTk9Ng2ppefGrt0gJa
jZioZUhWGj+SRaQFEnYMcuNC+M1jEHWclByC78dYMRcKfqw+zJN8KFzqxZgulNVq
fSK09LRRLyUrdSuNFsvbsT/xsY8YZD16kyt9KNtNbtOefMUqmD8Na3E1U/KjXCwP
qdJaoOPwBoJMKshUX+Xe51Q5uH2MoRagWiDxgKCEYL1q9lDs8QnQhTZ/0DY1IGNA
v2Cjb2SsSxl+DCrwFwsSgFMFYrhu0392aNx1cjVDPGOp3YrCCfhHbH7qfhX7YZmN
t863A2p178uk1BQr1R0OcEL1e0wFVpv6bTEawkYaF6/5hv+87+cKvMPlCrWqlDYj
tNSHR0Nv1uVKksIXo9a/l1WbTHJgtv8A/9FRb0nDtPSSiIOThqIO3zr6XbXrgYr7
4lqpmAOXfV5uAQ9eXYJhqLG7UHwfKxjmiMqVODx/Enk/0D56iZkOWvmv7C0TqOZr
iRyvjb+03ghtHLC9vB+v5Xe7gz8EogDeRpNSi0ZYO8FSy976gnJJ5YZvZIauZ7fi
tF07eBI4TYsocEbH+iBNaOrqoumiz5i22hfpJIrX84VDoWud76c1x9x+1new9Jg4
9czxqlOtht5FcDSehdP7CvQz2AV9bmICGCVxUFCtK8F8a9zFf6OOT9IxTKR+sfHc
skwHqTe9eNaQ+60/fOslWO/fHr+jeVJn9uUyhsc8RT6Blg1rJL9GCHMy5jpPHGaJ
qgAP/VAfzd1LonzlbFBpIzJRCwraly6UYiEO3Uo7Ydb96tHjK5zj39QJ0mmMyuNm
fhgh4iEU6aQSdo6QM8YS8Bf9c74E07/wtPWxowFW+vbXLYCQkwBxP4/RIJXau+wh
hVnqMA3jeggkdcJZ32zul3I5/v8cL+Cd52rVMvPHsMeJ8wO8Vc3D4DP4ciAge8Md
h4hykNPpQ20NZnxGrbXzIB0Nf4tAAVbNTvuu849QYwCcjrVdYxkEKTSt3uk/+4S1
O8dNBKmkH9rvjWvO4jqIfn1TEecyteIRmTubPD94JT6afuCKHSse20UZ1FJm96DN
f8Vpp8GgNlHfJgWQxdmXXsq5S/rRzsM+PK5EY391Znjh9oUl+ZoedLYxAwAOWX4g
FWIhJtkbMeJY4+Od43V11WYGpfXT/YR8PQH2oR8kc+FEgPdbdFm4w1yb6Qu75Gbn
A+1S1VvXZH/xdyWr8gkl3Hh/4+o5Kdm5cK4dy21okWDhGXlR3ly98PTzbh6eSlTF
41OvjrHtgTRcLaHanTgVUCysc7oXy5tABtHG1/NhlCsg4cpGGixknrZMfSums9LZ
uVATRORq0X0YoaqjMbR/zbmwhnHc8W8AnUiAttu2OJlzfToabjh1w8tJG9IoUz7v
7vpkTntXV2tCDd06RMTSyBGupl3Dd/Bg1XlmubM8cHnGKcEkyOGw6Yi0hhFz4guF
tSoV2gIJaJ18NJKkrZoJ0HxoxfRGFZiCDTEP8N/xtssgbe3HlzPBVsjG1Inwv6MR
N+shR943uGRmjAH0fkA9jTjnrVJRn1jO4xeCsGqbqGKG4G87FA5EZuWKAqXXgy+/
tnG7gxnjOhSBmQ351afZEVNed3D6IMU/9kAJKu3HAYzKXa9KGkcQMKzC7+ihM/a/
O/GwjNgfv2FiHB6YKQUgrFPF4+FUvwCIPZehfXo6u5KUgmZ1YPTYUhdX4RaSkHeV
eQo9hZk9rayz29KEzDjACWlac4fV0voN0HZ6Pweu5tqRY5vdxgqRQLRF0EJhgoqr
OFNDHpXFyBZ8SbO4hd8YAfbWbPObm3X4kPmcgmMVCgES3VnbOZKH1V9M2fm/WPvt
EPcTxfnxemxsACRNs7rQEOLWtH8Vxp/tLPfIlrtZPL6FNhaxvtD3+x8Bo0a+aIbt
sGv18r4BDxUggg5V5cahvMxpZKX06103sglq3Ss7VJgrbgaxwZQODebcV2MFWXI1
TRsnZe8Idwc/rB1kAleEwLrAOHbNvV3dcRWpueZTWKbUXlZgfg6I20KE1BvYHoyq
r3hwg40AKqsGG4wSsLwSiVHeHZiOCc+CxvfMjg2dAyBCxaNu2QT0uxxhhBbZIRVe
3+OYZEyJfItW42UVda9kvNR/Pl+FFiy5RZC65PJaNwTkCChHm+eWvz7ck7RHjJat
Qwahh1Pm/VD9mChG9EYFawQ/o+MLlWjuT0iNcfDHUnXpx5misoZbvkWZ1/sIEltB
rYUK7+zDB7DhlMbZLWbv7uOEbJn7CnaPJpdJ0c1ZZl/6zu68Rfs736laJeIPNFll
bPCXPAC1TtswKqUaGu6Pz6HQgsvBWxuvuOC9Ynbuu22TsjOaqlCfnMd23xMaLIpj
JhZP8/F+I5KHOuycYD9L/XdTB2Wafd3Sx1O8s3TFi9WtNdtpGqG06TKR0/db5WiK
qJhkpQq9UFmTnTIhb2XOr4J7XHt8kgacaglIeuU/8sNVCQqycTTAW2JHzoUf5EeL
g2lBIcpJCTWHjY4wv7+YVhQAQcnlNRbCgPna/yAR/+lVKxp7zupCWiLW97WrR0YF
6du6MP9hgTwFHtYM3TuPKYSQ6CPLHq1IHxkK1i/1E/q5gyl3LReZiM5eZi3so6SM
nl/L7s5MYj+fQpD/b42xx+V0ezH/fELrikONB4wNnCmFN3wxtK5Yic68Dop3Sevh
s9kvIem7okTPcjoA41j4MwLQLPg+G/zupEhZ+iwaT+MB4mPc4AqWn42mF2MfS+Xw
1aX6TJrSFI5YJw8j8jaSwN/mIb1LB0iOvWzY3WCeKAARpNVRtQHiDLipW/WAMaod
Dcl9tNw9uXPAlk12ZPapwVWx+lq6BosAGucOcuuXSwqhKhDR/Jm4MzMjVL7R1CXk
VpOtq0hZ+xWTIQTm5Q2dDhjmQL/n1GFiBTfunLkqtOAB+m1Fx0StdKyaIouIphFY
GTtNlT1vu70Tq2Ki9RORIaOznzBVEYORUz2gabyCos5rWAchop/kzrrz62nczzg7
hnet0M/+FmqrWbUfHJJ5iHKDrjJBEfJ/IwyJld7ime9zAtDx5YheQI0+dkiHXNO1
WbOiGiQcNN/MWGmiVUVGUzqZ4wFvWB3cLCaC+LnDaZVVs5LhefGxSBdUR1UCxUxz
8pKQmsO2CWxmO9lYmZfuLNT6E2495g4XZn4ywk4I7z4/uRQex4qwNftOC4mlwRIa
+8eRXOVEtvycvockJjVtrDarRANBuyFRsf25rt8antWKits+0WC+ErNbbN/QQNmg
08T19I/j7m5YeH/bhC9i+71gJTkvPVP/114n3IesVhezpzYGOlHA78uL34CBAzKY
bWUrcv72z4g0A53Ryq1U0HFukmpxh3fnAElEp9KcPhzMEBolJT5alnUOh++WnNwV
PbWVd1DjxRYJL8N/eBl1i+Uk/QRKXt6Fuc8GhzEXvZHCp9xqfPKClZhp86plNW+P
WwhRWETgDS3V/lgBjebGa9D1SU1UjksYB2W/vJQpPpCVhN/q3HSvM1lcYistIMKB
Om9K9yTNi1Y7ig8ClOVGiZtSpnORruYoMiFHCV8gZwLlbyoNlXKlQDVNNvvQxim6
ZPxYdoCf9Gqug0Qze7lqq/KlUKrYYlOFP+d90sd5ro7cxaH1XYfQTAuoqDnLEhH0
IcIYtLoVVHrqFLrQLvy2RLpziGzZrNVPpwv0jQM/zbMv5mfSIKbagjL3Ol/UoaF6
K7J0AEcoGOhpCi4VE7jxvY5wpFRaHhGUdrXQDUBk/pXiVbloXdixdQ4M8hokNUg9
hgEvGAKNamYmqLMG+pOiiSXzLvjRvTRlJvTadUoHNx/JtnhXXQ2J5Nb1wJ+YrJl9
Q011CpSgZLCbekvvVeUWM9252AJYY3ki6xNzt3OZZ8EpY/kp34PUp88i7o+ynLZS
1rolxed+47XXu3xifdQJ/K9nx87AXT8++cHrRgJLoygBP+XTrF8fXmgyEb7yDlKw
43kTYo+hmbDjR+t8e5gCFiuAa2FxCTZ1AxiO2eBHJHNvzYblTy+IoGzbUoBqrqiN
T3iqIr97MYslpecB7Mdi1uEXysQSezi8uT8XGaH39HjQL8C4HBqP5UrRUoSAacpM
lcyUPbtYPblcC8PnaZ4umgupiXG7RMrwjyBiajNA560DQQYSLlRVGPIJdgfnwLFq
Byk1qAw4NuZ1+w95rUK5zo5I5d1v0zOrtose4IMrAS42ku4WW6Crza/rbqPeGmJt
j8zvPjL+gQYZmodRUZNTyn9ASM/8j+KpwybndpMKzfrmBtL1fIDzT2L8NhbcAu9D
1EyTDIzfigvXXDLZ8+m/WTBGUwzERReBelCKS4gUn99g9Xl3+hEgW+1hit053sNw
FKhMHKbYlfG1yEmaHiWNyjraq4EwywzeYs75cCBKJzlVEPsZ6LqI9u6vX8AixrGr
xvSZFE4jd7cDXqsXAdPlRfBZ4Dz3wapEBG1A+NnUp79406kWzRlker9UOS6zpl9V
aPWUdVBoaPN+rb/BSKMkBBJrsCiMPzITgBhRIzT6rBxyUbBdtTYz0wD7GsXuWnGy
p0LVrge15PDoUf1ujE48pN8yg1jNjK9fyIMxUY+zYFtt6F9gHs9GUDCq+4jdT0nj
mSfH8KbZVJYibR8Qxt4nxVCzEjPHBH9pfuJ1A6uEWKXs3m7p5bgQXO7l5AkYr77W
oFFEAFlV0acErYk1wXSpTEbKIvSB+kFwxHtLjqwbqxOYLS4mPkQmBkGlL8rKIWj3
2K3s4P6v1eXDo8QxNpOuRFxdAWcc453hpN4Y8+O68hN+oaZKWbRdtUBt2e1meT/r
gVz/ym+LR8onBwivtmjuQEQ56TvEMnwFxzm0zbtZCODCy/OvO2mhCpYoY3huM6SJ
9d/3WexnbUajyovjZXh1TeI4nXUnMHJ66N2/m+pZiqCmWIPtfNdzhmE+qSZftLB/
iOU8qUnON0KgLf3H9d9uv8ChwYFpZXBFWOR4P4nKjkM6HHej5jM34K3CAGqRj/V1
L41OYwzuRtk1hKGUg7OPmqHiKnsuuR6Uo0eYD4zfGUrYQWUKP83LtcHvOcU+o8Qo
yrtMhe0nvfptvNy8aZG/s7C/7Y8QidWIqob4ZtNe34ILLcO5IOFdb8R1D6TSFmSU
NTEq9tix1uRfOm4ASal84jMP1R7Yj+JiB9GeqsldYuBWCsKQxqYOsCa5Hju/l5uo
X/PTX2SUth696qFui45zLSajxIwNvpZUOHhyIDLq9tmxhglfYiC8qST8gmiwzqHv
bvn4wxh5nockWrhN3RDyOtFBYc7CRyirnU1Ox0K2W5kzcY9zVIMF71n6fK2e1pH5
rHuTsiUubGp2e6Uskr6xSD1AyPiPTsHcYCJZ7H7AcduA/q2moZgdywDFv6Wn6IVA
KtvbO6lIrNBNyRSn4kLfCH5bVuSGNHVNEs1LpNL3mP+1/FOemTK+xLiHlfDaz7wa
QXCwtWxoCJesaki+CRpFWnigFmfGA9/RAXOOwDKutIQKhShYWZqSpjqBD/wMoHwO
kxxcnJiPO0P1DZ8TOrjeAphdMfMt626nsXBypd8FMrSk39keiXpbe8R5rFpK2WqE
/7A3fJ14hJSkRiYfEXSWTKJXAB8MbDSmhp7522TpPRcrU3a8Wi7Kt4cVVATuyMbr
rI3cviJNg7sMmGmuhmXxjRbby1hcPeCUHJrYhLJxKA+BBtfyYoUAfUcwi1bsNOiv
ggXVqKM3/ZdvFhrCnBSyVNO8k3Hg0Divc85Ik2GV+Gq1xFo1syEyzor1WvKzj741
z1ydx6r8XenYW9IuUFlTQR7aMjs4QAJlOH0y/u5pP64aRJTVeTBty1lCw9D337PL
xmgvO2APAhMmPg3gb49vJpR9S1LA/ODM+RMAT6vGLGN1rMjPvCRJMVIZUbZQPVBA
vvDGaVS+xM2iLfuX76aZSuBpMO5ODf96l1PCU62g/i4//Emg6wsPrNrr1m4Pev4j
yP17tNKcqe4e5sOjCYLeyjrOW6+Wwpd3W6yGJyd+Y9OEjNpE0iRQyKRAfawlrdpU
8+ynRGoTlX3K/o/bnbTR3b7OavXJb9wO2qHQkbHMQKq/vu0c9mC+A9pT2PR/GqAl
V1AJOARC5FUnGgneOVU0z2gaiowduPI8J9tnpIcBe5NiDXmAmH9utQ8QPX5i9kpl
wVlbPfewCWbBwq2IDZI5ywLgy4kxph8U7oevx3Q43Te+d2NOlexMQlxvITXK9hrh
MaKLnP/Tjc8wHLHTWgw+7gBPDQQT0Tw+N5wZuHg+IgG76it3tV0KB62n6KlzNuNi
52w5YLZaxe43B58DYP1tAft27GRiUgwMJxj8UfmB7rX0AcBFNcKlEaI59OVu2xF8
NfqFXkGoYtuyps2eSL/MrzfqGgkl6uDFb0IZjX1hoXAD3VxOCC/a7EQTJrIhJe/r
YgYMF3RursSOhCqH+GJHlaLHtCiOBlS7Q1WFBJ6P32r0orm0wZKFzAOjFAiEN6JL
1ufHOaiNNPleXT2VHZ+LByCSPICKKzrEwcoSjneNmEvKOA8jhNGekK0TXdi5YPPQ
Bs/OWzgja5/wqVCA776DHdaX4QQfkLeEUL4nroMl3QiK8lA4vaAvkHw/E8razZbF
Hp5rBVxcWyFFIwuw7s0UDrF8R1aQGnwp4ehhLd/vnIcPwTmsN/fHkyyMKCDnSAJ9
i12aPb4NLVUKXmc5C/cy0K/g2sb6KWemyGetexWr3c6f0E1yqyG6Cv7APRAl47sf
M4QSInhVTMY13iNTgjBm6YTVUAG5ggi3V8vhN+1oSRXGaujJ6HVzziw7USEA+k5s
/XccIeV7W7xzzZALaY2Tw1CAXUWMM6+UCKRFICCj1Yw2uYCLCn5CUTrMuVwfLfc6
Ll7/pv4ZKrIYGrkBrE+qN8hOu/6l+6zW4W7ZkP9KeBNCaQ7ELxhtAOR9/12n44cC
h5WJf+HrMtyLe8fn1eAGKP/w0j/qQG36J+uLlQ2lkhFZypcEb+JfBMvyWiSn0e5e
SNDcQmtfnN6xw7SKbUNZCnyrip8J2aTMJgeJ5ujw9DUuoC2RAhDPHpbX02Cn2O3j
i3hPxUghfee80SYRfO+AT+EYmb7DC0mxZyb3AzkU7CHdUpEPMlfGZn9CIOcTVifN
Nc0zrVZaLiHln8oTxpPPSWnHU+/5XEl+NEGiVEw9Mb1wpFbJSlkyFgbdot22xGd+
+ZJ2ippU4bVwJzthdcw3xDe7e7uqSY/KFb+CuLtZOjSwo/5dquGJdTdBfIqAW7xz
6a2MdMLC/25AfqTuJgBmjX/C/FYnCfb+3hz0ak7dxh6CEBDGlhsejSgzDWa7n8wO
dUs8ltIil8Jyb94dP5EBfN/DCkULKqyrSXxJ9uZSd3WxUA9uBxoBksopF/dmzFF1
+KiHE0D65bzwv+TtMcWIZ8jGXEPzzCf4wg9Nz1hon6IwoHPfqDU9AM/H71TMhkvZ
csKqP9ag3tA1rCCJB2ifQG1hCx+nQaq2859YYhoFfDRzvokghFgZUCsgS7FJjhlp
21cjy6EgC5LhrVUGv6huU1/3WatkTNoGChlbg9bq/nEFqBHvtvKsrPEV7EANoS9T
E5z1ikojNSI2HsI0KC6xRNVuv7dRefWzI26Z2OP7/692TB3cO+TyeLvNm+gtClT8
TaRK+AVOOwDOoNak8zDZKY5kfHj7HxzcowdVG5CgeJm28y9ZPGsKpw5IaYUGBdSK
y1wL7yn0zkzE3vHr8K51LHWKxgznKa6F/FThAI28STf7QqqqDBdZfu/iWEOCmmEN
w7skoEHF8F9TBaKwHbFJj7EKEXZ8u2Cyr9CYygq7q8xONQcG1lqQxERaJHH64Wwp
1e27j8Om+JzgUdrMCg9X51lFJc8gVgWQVwc5lJVfE7rczeP8IIynOcNtrlG91aIx
o1TWdUzA6UgfjUdAP4c+259z3sL5QdzvHoS7rEvFtbcNJNy1pzxWhCh2WRbgMbo0
jHsSLR3FvFqHX05YZPlstViBb5wb71Lr/jgP/n+lWPrpkLg9ym7uhnlDbYrVwp2U
ciB5/Mf4tuN99au+23W5kSszi3r8XsD/NP65L/Sh5LG7RnukeL5xRvrUDyVevRLF
MNlSwVlnaYqY/xQKwzMRv+PfUHsM5NZ0hWnpw63tny0vCEW6aGl84KW0AKE+ZtGM
uRa2DyaOEnbiNROwUTGHPX9kk+iPOTSmRfFj0RRhH37CBXQuTMtM/IVqGBgkGNhT
wKNkYt4oF/9+WwDheCAuwB1APraK4B1lqO9o2a/6ZVz7E3lCW82ZPG4vVE+rciV0
g9t76c07mvXd94U6gHp1KiVjVWGcNNcIAODhsqH+6j2DhXgT4CryYSQiPn+wXg8D
zrYEXYJfCd1QaKVe3VdLaFGsS4FJ4+t7MS/zRt+tjjEPDvXk33pQhoofLfhVD9F6
ZZqbJ4G525PdklHz1TkohiDeTomKkmNPcPkNrq8W5lV84Sf9kbblumEC8TL01FdP
6HkXb2C9bP5UpMEPe3UzDXthu0zcfmPobxHsSfwCYf4jIAHWxXMA+7J0tvtJ+SOg
rQdo2gN+WDBt9USYtwMbX6DQ6mzY24wAWBKkdZYLkcm+FX/NjUOVWlIUN4DZXa0q
vxJPvyOTsMjAu5JVQQ3gMv9EBl0X/qDVRC95//9/SNfe7Kp5zm7oZDi2RzH/CD+e
2zhE+g/w/cLnesFf43yPJ51Qmu15WMcVhCuzUKllZMgJdVmUocxtZ22derE81Zn2
kEJJIKVarXR1qBzfPzMvj+BUPG84fGu//uP3nzbq774BC0ddnqTUAvTMhk77M5w+
C/uaFEg1RZFaJQ6rDRyFUuQeXtzqmkHk8vet4jydQsysA/AcUVVG7eBwcutDK3Dd
atFrBY2AuyWFM1lsU0qKguWi/FVs+3Mn70SY88pq3KXxcIGJxv8xWHQXw3gGrz6s
N+KEmzp9QH8+XiXjawx8/Gec9NvhkW4QIF53gTxn6ZzzNkj/lYW9Ge9CGtxH4ft9
t9ddn2ytXywaHYYJRS9C+7nZesCiS1AwtPCTfExrh27bqAlIWvKBh7fmjaXWQLzS
utfrJsfT6hdDdyIRvXhXTS3bV2MaVGyBi1qKKDAl7zozMwM5Y4ka0SHCee48uX31
bkEB9L8201V2i3fTdiwan/Uv9PPXO8lzIxPr9/VtdTawfPDmgiufuLYJbdOFLJnY
LQBYbTDazg/vEhbaRfl7/TurvnQeDF3Ep7nFSrnEeL5Mog0UA1Gj10EdSMwMPqXs
Qo98+T54/xuz5LHtqZ6bnRxjMY92H/D39h0jtZv94Hx+ih04GgANgS8XgIhM7m7d
otfYHfFgMRG5AFkSH+NzYSpqZaCjC19Vgyf24FaHrw2O0MTRa0WKGmvmi0jKneWw
H4Sin/DnRGEm7ksmE8FGHg1KxhuTidtWA0QuSacT2xXcCnUuDha4eprRRNBpAO2S
48/u1LAEJC2IlYjVt69XjjZz8xfA+llot0EtKnUt3M+uquBUY/MDKyyqs9jlMwvY
T3Pz0QOHh7vMR8ZTGJISziy688f2Aj7dMUyiDDg0ITkET911/ly7qsFEHfhY+3/G
idWm0+EL9L4rUDykBuBC68Ungz9mLVwWTcaFxKYSbcIyyaPeE7rz12U1sAVGD7xd
V3i40HYKkR2tA2UCygOoPgVGy+zIgnC/63FFFXg93UNucKOmCNlS8sGTDqKfBSQ4
W6YRMIuIO4aM1TL/mlwrmyyngYSJkqU8kUnhbWGMC98o17W8wz6j/bmBK5IN7WAi
ZjcZQxXL5TuGi096NnZoZVEGLKjRUBbo7Q7qTHTwlnMc5dIkRw7y5sRMTzPvaZkl
IGG0CiocCii6U+ehXvdowZoDi/Zx1I5VqKEdMchfmj8NxDdq4QrWAoHwa55ZluNH
ym4AQDPJjjZU4mcjhyOcCy9p7HttOQ7wzTDOrKUKuXlWiJC5tI9FhiFice53RVs6
+d6ZhCLR3Fi1s6NqwwzzI/cNv2upTB1r0k0o/mW5X3Rgi9ZwO/bXaw6r4OeaAYHg
NiSsjtua1iZht1FzNXmeBKxsopXEqcLhLgqhG+BZAlsEPsYpSj0jWzuodcDeHqSi
SOTUD1cCitVyYLPwFYy/bT9lHpskyi6c0l2O85Ef5dVSw1bY6MIrYI/cL6V5EMgG
+vhRw6F6quaU8ANIqgNM5uOxyab1wG8l17EekzWia+W5kT/fW8XLYAU0z28fjT9a
SN436NmOBjDzeeZEN2DoxfKwvwGMH0hipRLR5zFHCqF9T3ki3yD17b+xiFiYdZLt
I9v5jniRhP0at6gEabT6BILopmgDU4nmT3qEWT/i5ntovSV7D4wKBY+phNfopLkU
QUSWofkEUotr9ehKQaD0YYdNfUK2jr2zEd3kE14ptzYtHiQ2tyBNU0ryAlIO5OoR
FplsJ1vCJnAJ8p5Q262nxhMXPYPINbevAzB3FolpodtpF5d3bpQ2t807yIlnStw6
NoPeeixQf107zvXEH28wmCr98x8xh07HIZSi8Orxw7sH4O0wKijNQv2v+1/eNDCi
SJcrk4X4Ple05QuxpzhIXVSFm8hqciXubBXJ0Q62O1iDG9UnlFA/GuNefeuHW0l2
B9gTnKLvyHyaVo+PgjIePrXh4IfNF7N2HFcm125Wv3NdDAfL1qYd0SowdIcRUDqu
yqhlRIJrLsgqANUhXzFMiL0FhibISUPVShv5kKXdkjHJrIAMIXrKCciCOfObkEkJ
TdZuAJ+0QRyfV3H6va7e44KOSGk33xEu5tw5qDXSz30K/LT4eJYxKX5LmLGgVIM+
OltraVUeltLKChDtSd9Hhkw8cJVn5QvNad6E8j5y/+1r0G8NIgO/lSa//5ukcUHu
izPOSZrdX+lr3gAqsXYVWc2MMPA/ewd+tVSTRYnNjAvgJr7sQS0RHc7CtTyYUnGM
+VJfDCJV3GviEVXk9u7g/elwiit0j9dHp1itu4HwEurtXtBlBwofprErgW8oGEu0
2wHsoa4SVrV6vzJjKHx6YByrqG8e0+3+c1EHBWZ8+Hcl5ZMTptbl1QWK9C+IU5yU
GCFUX3OR0UQOt85SYgBJhrCqoUmyxTrnXGFYSTsqK2fAqg9CabV+OcEZCF87a27Y
PXFq4fZLzdyyMRsupzx8vo9t+Oh9txF9ShUpv2Dbc9P6HTW6AESMPnVUx/OLCInJ
4uhEc1yPXTxYK7eOOrq+f9TSDpsPWLpZuUGeEdwfxS02628HIL4yGpuByO84xPXu
jXyMZYFimufpAKJikFJrQv/XCnn1SjhOtfq+y8UO8LGJ2n0qqFGoYusfNVsvosKX
Yc4GgJreJDcP6MR7nYi7SzbGcd+cE/Haubk6GKERLRIJYHOkli7INLm/8ClPaj3W
+CC5vn1BZuyviziCumo3SnyrQZTzia56/QtnG5A4j+RMp2Kml/ZW7GIN1NKfIpT0
aIdN3H3xUqE4FRDpGZEFWdELfhYSKOYFXrB+2IjqbP1vX7UG1AOZre9mhqZ4BsUz
KcVrPsNiJxmXY93Avw2RfPCdO/fYsgpdjUgvgzf4YJFjCcyWyT5B/W8HTMckG4IF
HxmyXkigiyNqdMWoiSg0QMrkr6z8k47tfZkqVM4kHvSfskCk2KdFmErTQJ38AvkC
YmoG77Hpr6TmbCdwE/OhBsG3jH9ISuLw4hI/Cq6X8XzXIGEgED6ikPiYaMoVf6DD
8GNiefbDaHmel2cIFhYvANUYWyMgrSdrwq2jnBYa/FgeRjzmOEYg7IRnDiXuDBwy
l+zSGeT3jueF6ysOPw3eC5TZ9W2WFQpzfgczaIaxXq0u475wPEfBzDYdO3xBUr7l
zrippvU1Al9ArCXmiWomWgoruTamPdWH15BSKxDwVvfSkoUWtJreLGMC6L9KFbh7
XAeh4AIP+hJl+68sHX42xwAsUy88tYIZm4L3zP/91xn0xiJce1FYW+utH7yUjZW2
8ubrCuH48j4lPihp4s/OmWRjt7q+8V/Fxi1tT3tB8SCs9joNO5Y0A9IRQ7qmXS1d
oIJKev2roFIsyht2SvzUWocTW0RQAQVs3jJq3cLKjaeL25q/QCObO3f8Ufqz5w7p
P8ryze+d9LIkW1nv+vWJ1QCGrBPLzn9jaYqEyhxyt9GGOHg33IHxLs3TL9ML63HW
EKYEkTelUddqKhU1FNh/RpjKcW1QqWZucmCrEBz2THCGALzOeYTnVLyS9+BQWGKG
vnIh6YhNBeq0hn/IHZ8a0E5lJXN8dzH7wxep51iIWy+HMtCNJog2RoJn/yJ27ZOx
MnwEag1QlbbQ0rq8qVS3FDJOGWHFXzgy/n8O40guvXI8xOvPSuA7xOxxQkdXBRDK
MhOtrdEeTDLxk1Z329nkBYD81l8SdDnEPBkwV7rdMmEnF7b3KM2R2fGJmAcEvQ2h
84Eh8xttTQwVpDteHWxgn7iV2YR+vGEXvxHAKRjc2vmeyB3+TU1BzjLvsTBhwGEG
6XGE+UwFXKdGDhXV2ebbn74RSxaRpAjveqtAW0ytyOGYwXekmSJVRlzrdi/IGb4j
lzUa1Jd9yrHuferZ1fgiThpgOn2nZ8R15tdEa2rakfm7dFUZ8ah9ZcbYp0BwrU1F
5mI+ciu8UIxjMGgL/zuDEPIoatywAIvtT7oCxdxmRheVBhwBodXjY/ca7wCltIh3
RZLUocGVUx86LfweL0CIvLgWNxAkm9mv6HNgmapOqak4Q0AuQNZmc6Il/XFYRcBm
a/L/+x/mOe9I/RHpagcKCtXL3UI5bdk+5MTE8tP4tg6XiCuLxXevRli3hHJ/gGrn
6CCMUt+XVO+IM8gFpUGEhHn7C2y/0AG2+9k39m6dbIiilezbb+3wC5v3PXdWKgnA
vZnHDQU8UOPUxki4Y1Bb2MPEXLYYi2K4nGJda3galrbvj9nvWPaij/egMusUAUbo
U27A753Ctto1pSr0Igh2Fy7VfqHq7I/W9EdWowhXQcvlUYkD2Yj8jb+rHZvsXJPT
B64JBE41kcSr3IQoAYpOekal0fItOXoXaFh1S9XDVsqfccJ3UdseztGoG5my5fGh
ta5XsqgY4IU9AM8IyOxUlbtaaVXX/0EavwPwU9kuHguJqCnyzaxcu79y2Z8IMDuk
JsaHs86w7p2UWex1FvVFN3vf/f+FjJp6Fx7SER0wGKMez80q3KJM6jhn4CnVXix5
f/oKxQqhRiA/vgugo5M4NUR03PpURPV9FpxMvJXBoOHZnGiETczbez4g7UUSoNir
d925E1vJ6KHzwAmodCqHdbyK8r0uXObA6qKjXDBmMgenoSoZ2ClFC5qpKknn1B2b
51U9p82Y0iu/0qLC+H8NKLyOij3yBMWoLA4ibhuOVdSSZfwrtAWQq0TasJ8E643A
7u94Ur50FjksrBSl11s+kWKzKtRUtsVtSj+i0p1W1lq4675dOZFhk0hOl9bMcvwv
zjMlb6PLi6cuFLyLsP3I1D0G3jJz2ZfS6OxlbWXH3FCsGGa+JuytBErGhlPF99dh
AgJy2AsQQk6Yew8l7rGIJ5fDUrRT5by/E5yaaVvj9oupFpiL+NmCSCGnACgOgAsF
I/tSjfYwlSKmvWP5dIXGZwQlUCGcCZKK2KqnRT48e1a531jNJ5B6b/YWEtcQ9Vfu
yN/ktNMHYK8XlRZHFTYf3FLzNYJ6NCQJKca21GbKblxKTitZVAq5S+D9aUPt4dq6
Or4XqTx0PhuvlnjTHAMKI5Mk7B7nBdfnVJxUpJaZ0mBpkH2lhCgsbok4P/oyFO4K
6OGbvfJUkO7D80QfHY1CIrvT8u/gTC5kc576mJ9fnUqwsb2ZWsmKyPxGiw7zvaYb
ADbTeJHAWQDlZSymvFDbBdS/lZT+TdwFN8Yr9NSFZCCGy/uxOwbB0JRgb/Oi6gP3
EPbQyvSxpM7OxcoqnAu8FRg76iDg1ZYZgdLyjGClCmgYt+Mc2ZfyyA4KtsNtca2+
o0/T0GFVG9gNjf0wnX5z2quzc38DX8xyP1T8Lc4GArUPkTlk1U+yQVtECMgnlDc8
+YnfZVziX/fjcZMUNyRkRnXgymuJkfF4e/iEIyV+fPedWXpwUb+iS5jEwCWMhfCx
km6PZb4B5cls/abu86k3jPzSzTU32RPqtzapsfLn0tmUWJikuZTz4YUQ/QuFN+JI
jjr44zz4SHIhId6dlJP5VOE1G2BNjwGFIvyC2SjyvDurYqBSs8zWxBbsqOkGfPkI
cPO1SsogpK8xnXZLqSoXIGKao3AB8GjnuQ5wcqOWkJptPlNjLv19vmLSoUqRNesZ
dm2lXKp7kqU5NgOjTHnidf7yqYijSKE5wB8hL2jrh/k3E5Mrd7tprEIAGYFvFoe7
3J5zg6AzF9wIiS2p3uIEmo6vBPNw/r2NG0ahEdBF3TV82aBabKjzPTPlHhkwskYQ
AW6J3iW7RGr07UKYIKCqEDwQfZ9R8lEX2G1w3NCeU/8Nqw8dtfj9Kyv1ZSxA/Xs7
W0d8p1QzelPYqTfNSepv72WRM0x0THIEcOvwD9u8gWdG60LUswoWAB5jWoyJyNAE
GJKGiqttIQYVDXj9QrvM1bGO1mf3GvUxhJjEmFEeizGCN4lj0UzSpHiIVX2gyHbX
7TWc3RhJoUEyPAn89utCqU/kAmFtf0TUBM0yT+hbXu5ATTpvfOxHA6eOJIb7Ndl5
wOXrm36sNuxAxGmvhDnDlLq7MRjJL89SZj0xlT3NdGvMD2E0e7dHws3RJM5PGfRV
eL+IrzGRo4DKMREMgYVHfs/1FnkXbaR+Ksz0nAe6MYmu3I4LXicj4cS/tWJKCOqS
/txxprVgpWFoHxut9mjvs795WZlR1zk1l6OuHBpw1khb2YGFcDcSV0UVE+X+locc
6bAdC23zW01rg9Ivcw+ZYxP7JTvPy9a4GFnwKhpQQnbYmSCuD1zzvYuIxD4KCJK3
u463TETza/0Roz2aqcuFbBwNxtHchB9evdG978RVdafrPv1S2nmlAKZIajU1JUy2
3sF8FxQ9bB9LvV6cxwA/tzL42HHz7uZ54HDWOKUozstj7Gl1BT29RnwTV4lXIhA3
rE/1k5ss8k/EAdY5JPciMX8FN2go5UVYcxiNDB4wErymud60BtJgNErVDmiekT0f
onvnyzWJcyVeRR6jcEAP9Ucb87asl9Bv1s9cTU0EI9+AauU6vmJao5j/30UHORmS
6Fw2D7RNmSquVfa6A7OVaKoiP4QpEGv+EkzPZhaAUUZLiOI8oiGVDGWwcusU215R
1KVjHBjHdukOrjqEau6EULvIiVXohxKIa5CRNvj1sQshjLv2LVBtRV/APnXnmai1
Ci6+dNg1B7/P0NyOcsaaod2go2JWR304v0yTru1PJkNm839rvP7h++GJTFxqbkD3
RbT4FDzf5EGjGJnDrE1BzD+9ifuwbk+rI+YFQdJm9hDlF9Py9ntMW9/mjoU+3Eh+
3oHKZ4ypIoF0eIx3mGvjdbFOUnBkPCa9CuWYjbfiW6W6k+8kPEbhgBSRF3nUgRaj
qXbKZncr4nsMR7+gQa+NbccL3f5icmnNiklAcmt4bmPAwgOtS2G+sPHEkLAe6SJv
CzKa2qQT7NLeM4MRZnILlsAfceePOOOReQ0eEwTXoA9fdB/RwNRE2PNpFjueGpGg
X1/AX6IV2sQw0FaJmASgzqfT4FgapmTPRMTDgPA0vkhE5SGTfyykI7DjRS6/p9Fo
UHVPbKX+sobxt4TyYOFQZvZpVN0a2fq0esiJ3VsgoM0FGcNreDu+9w6y2tCejS2h
VlUqGel12yUC5JppiUIu08PCNOE+mfrZVFVvMInsTCly5zCZjMj/ezZ9ZHEQJi1J
xOoOIq8obgql/e7tN2SsGf1MCEbPGV4Ia9UuLSTbCRnOXDCQSos/VFsjJZGgbCj5
/Qm5V2lEAu6cV2UQHl/uhprE7OfCf399M+Ffspa6nrogIejvrLOlR2f1vMeHDp7/
D+dz3iSNB1fQR/HdaEumf1Kl/fjLNwInPuxYLCq05Gktw1+nqonrfBCA1HDlVkZC
4DZduK4JNbJD++x+/QabWnjckWypgZc9LJ8TQhr8O3v/E/vSoguPBo6KThyqcBw6
i/vO83e0LXSSVGxC7ANEHM2H2pa7HZNhezyBQG9o5MGrOKCUs6eJEmRx0m40/nhQ
RG39miuyRBKnSBgL+0Tm9NNcUviY3BvNJPwaqd01R4fZVKwAvRYP4Bo+btCrwapC
HVZpEcMuOroNfWqss8Gs9sgqciK0QWnHum/UDT/c3DF9RlQzYiAq8XoYXmDXeu0F
asVYECVQ2vSt0MRUi70vyV5puYt6bIacwnOoZA4dlqfV9TBlLEYWU43rYzPHlSqF
p/5FnmFxD18czdgNUMrfuGbwpXBKCFDh+o9t9BFG9Q2ZCDeuTpqRZnygviIyoSif
q8ZXg7BT6gngVK3D5Ip+EGBWuqwwp7DSlI1cwXRlFPbEXZT0/ACzjAV5+uavmTo6
XxWf2DaldvzZ6l0Phtdg9zWbK4cc+iaLhhj8J/cyJTXp63uE9HcAjGkp/34WQXkC
j2YF+BkWCHTEuIutKHAJ1zrrMNZB6mN+dJdA3qGhuG/H77ivsSk0H5DMbwyh4pXO
2OSwiHlKKXrUUXp4T+ViznoDbJMR/Lom2wNVzxtSHVUPbHlYx1tZmolO04hawP6K
6AVHMazBHhY3wwmSJY75WbGOUufwsK8FVaCOOVQaaxuHkDq5cvvmOVqTmbHw+ajJ
YNmJh0JX4Zj65Al1AbB34niWpZxNvd8RWDjbhxCgOPYHjLcl+Y26cz4KL8DSDZ4a
cNuhlGQTIwKuWWKFKVYTosORYCrk4He8QlwrRDJ8XJ0P2Efw78E8d2m4ZPfcd/L1
vSjriRQFFsU5IhLnng3P3P3t6ZisdPu/g3Lt5cGCb4G7kq+jWAOIml6ioYU0j5fS
xMtuO7o9nUq2Po6udaMQnkgdGx1s6b/bECcSO1H00zcGvu8aq7Fjlq2q4bE/wbA/
87f7xCoVTlvKxx1HN7Ju+Q761GyRB3FuVm5VPMP3MFFvmS6MHmvyk6rM4k/KWTnI
rG5NljgZ2ofVbtKnj7QxYZRfjaE6CMGQx5AlvAq4aImWNNLpV0gDOO6JGARmFqrD
oWGD8fxlMvgCkNbyh52Yr19UIQZeafYGXtCFv+jDk+1WRjy802f9kDLkDqwmMBlt
A3Dxy+JyQAc2xFJ4Hufhf/IvWsEpQpO3Q9tcIuIwDSJvtDXPEbTQlid7hPI0vY7h
iz8S5VYCaBKH8w8o0P3QZboWCpdQh/dHyh7GN16IZpa5HMZvyCL7w8MOweCrpRPd
vDdcLCOm6D1qZAH7l7oey6Ldwaqy0xGGPw8L+Orod8dqymQC4009iY4ZoVxngX+z
WRju4XHSPT0+4mwL63Ht+LhKPh5NImoQWT/UXzjPWDbkPXwWgsnQ9Jgcrkm3CH+D
L5ehUR52QwFUISqkmQaHAATPnzWiNZWnci5Mr/27d/4Cbr174xozWaAlgDL1t/zY
Kuq8nrpYL1SGDmr3hHtuxFe3rqfb/4CWdDJasIpWvRpN5yBf1q74rcRoAgMAKWo+
5X2MEqri2oaQ4PTGj72+EsCx7hza6kXwsQNTvQxnjQJqEBf3udl0I35OmHBFCd8N
rZcW6IDvvOEYwK1So2n+BG8YZ9YI4XHcM8/TEBMVuu6l5JmizuybbBiRaGwoiLme
7hdLpYnBvanef5dgBaOBC/LQfNrx0Qv3bNOE5SnMv411FPjWgxj9+MO910/k0cvv
XK2v0jpm3yqKttjmOuTfRf34KLE2v/vczhKkB5O2zIzqaskjt0FVrGS2GWmd7On2
Pud4bDa2KkQtAznoc83iYwmUoyOkoLhgYToZPicwl5Y8vTl/BIp0ufHB18ugp7R/
dbqgx2MxoKzFyzb3NbJxkYFaAgI5ICItTgdPR1STj3W6l63IdUkyArtWq/mFejKS
gh0TvxH4G0HTeyh6VoYwIU+Kk2y84OnH71vqJ6OYn15FT1Qcoa2IvADYjN4NJ39I
8zn0ljgIq7pyII78RKwx0aGdD4HJKUZoKBVep6wVL73CcFDOugWw3qlO96Wghpv9
BiIj/QMLpBQ+sCNoN5DoGTaqdMXlMGzkfusHuneLnhvqV+IsEP1uvyUcDcbJeP3E
6TXPmZ52rBEJAOcqz79LUqpq80T97bXVHMIHCJetq9o7Dh+LCF798VsZoRsm/DeF
WX9/LaPCKCPnHLulOUXzECM2x8ETJaOc9VnQQBnDiXCtcDcBNEH22P4W7APVKtu3
boTV9YVYTti5gvQzbYdSrEYxs+iN6yRwVLKDL/56Z+SG7IazMoXkob5J0ah1o4N5
NbG5HaRvsBpDKqXEub/uhJVlKCThPzwJwfxKdvfr35i2ZI3vohMYr3sdzJkyFZJh
5vrEWPKySCiaXZ5B8GzBteGp/PyB9TgFZwBrXiqrQL4nfDVlc0iGzHWeflBufVzp
oCwFRMaw6mpj4EceoShiwnLUQVQ9Ck/C6vTHzWRBL0rMRT7k25EiNq3yBzNcW8d9
jOs6HTIgxaCKBY37i2PEd3N3oOOAWOkPZk/xTfjH2zeOVgO3Utt4GlrbdYajd88x
YIBR7WXX+tHAwhJe6Bx/o3ZqD/6H8N3TT+75WnR7nqJZqEN4zyncm/JlpQW1CbHV
V22lSuMNiG4amBn8WkUQKX8YQikMd4OVvk6uk37xiN3ULHy6MqKA+JByCMmubGSF
xtfAFISC1eUw5C4/3HtqkQUGSdQtKVSeSa15QHVoRrjzfPWPMh29gDE5q5AAihXJ
HNTfHdudxB7deCSAkZ4itskrelQB1SFZyqCssEQy/on1oKVLBgrsZo3HZ8+B6OQ4
su22G0NdQuMZz/ArUgQDcRwBoG1vNgnuj2vM9TCUhzzVQkLgeRxFh+TKsF/6tRcO
0LgxzZVg+pp3N/N1n91qIKIe6tu5/vZ9m+zWTuQRf42mIkagYJ2KhRGTzeZtupbM
cPTS9Y7yk2xdgMSlJJpQns61OxzRMXDHHjHD0xELPmDqPtuZ0vNz6UQBfSBDO8Ms
eBHd+/id9qEp3j7ecuGgYp7QWNhgtTmGVTrWJVcSEMLc7CrKCwNl1pmkGE0Kcb42
eD2ZZztW+w0yY5t7YchzN/I5DLari4XMyDLc+r/GKhZ3ABtBH1gttxX/59weGxNy
IliUnNXUz4ogzgqKH0mBDEaCaDOm3gU0VAO2hgSJjeY061r4Xx1uaaa8OkVI/Je+
XWWoYAHpUoS/phWT+k+mYePw5f3Ti5RsvPTYmynrO0Y3i7yppl//jK9JJGwLMjKX
Tz+hwxN5KEJNNSoUd0S5jOvl4FSJDh86rGv6v6evkISYixJuBZJvoH4XS8DK/NkD
QnLx6d4nbnyOfkkw/ejhG+IgCWln3NUEvVroI4xBtz0740rBF83FYV1I/sal7X1Q
SX5Sw2d4gpv3Ftft3PLinkkEwveGQ2Mvc8Zeh05px1DVq0cdK8K6mLevZV9YMKMZ
M49gkE86pAji5f4ziPLGV2u7ZgT670+qpmSRRibkZ/FeFqHOaKVGd/9ph44pqqly
TVhj9UGzDi9BIiFR7K1pP9T1ZRGWv7pHkRAGnTzy6tYwZV/cj8qLcVBaGAD+aOOZ
tiyg1PPPZ0aQoCDjORjUStQF4cntQ3HJkRQ9z4NQ3n+lHyjQHxLbsV4MyF/j88N4
wnsmb7J+g8hR5ODBfg8OOS3UTe4op02aSyC5QVBndfmDDhVBHzon18Bi6MovlxYb
7D/HIGhHU1wlTqS1v5/CKDKRjpMZ1IQ4FbDhiIkGafkM2mgOsAvzRwvG6A6Q5pP5
QKKcD+bJNTuPiGePYOjv5u1iOiWFMIsMsMjJjQMy6S9FTUDHzWnlUlCoON4v3Rst
96hEF5bFtx4MGgt9TH2HszbH7C5HULgGaFlgcDE1+wf0G5RUhXGHc4Flv6Hrl7h+
y2NRIQssEQZ65HvAmhOgDiyYc1DiMqKC0yar0j11mPh+himCXoBwiCPdntAoeVwJ
TCSNjvx6536hXhi/eVA5FwUlCQmtsztTxEv27gLwTBhKY/XYEgztzia5d5Pe0wU8
AhN4KE0JHW8PSE09mc1qVcHApswPCjVAR0cQ9aSjIuwVGHzFJDx8vnLqLGjLXxqY
ESQ91RILMYFeb8M1xvVgI0gdjZ58QlzfHp057gWMw+fLDVMfx3oRauuvLQDICUpN
V0PosdVEeFKSNYml1ULWuJV1MZJONXO3GtFBtfMBH5eXXmPS0qJezG37znBzfDHY
ElTf7u2XFOL3xEISHxtATzrcFtfy/lF2rogkSkf0wwywX2r33RtHPWs16hlQxqU7
AIuF9W9KtNMZS5qUhyzsqSxp35JnbRtUBXzm4slFMKJNIkYqHV00r5mnXxPjRHvn
WTqmGAekg1JRCgJ4JnVBpX+46upV6oMidwWnTeTHC3cJbmM0oMv6bBgSDBWpLmRQ
lTVQA6TCODuW1UAbcVJmeyxqAehBzlQOeonI3v990v/PpAEjp6GXUTK5QO+WvRZN
zWOup2jsv3x+YhIohujdcIEzp5RSyjETT45ExRgB69P1u+AUDtwhyYVy4a7V4fuu
kdLV5lRC5wH0wO0D4gqRqNaM7ksB3OvK0a53Xk6PQbaxkWxZCB74UdfjXb/l/4zQ
PapUpqcEXoDs5YnvvB6vp4qhCMSfvsAtogE6NNtukio1cBb2W8KQiQnbm2T0Be2/
CleQACmsB+lWLE9WZ+1yf6hdh3KeGRzplaoUw0s5OHVLJATFD80vRfe19iCQodSO
fK+G5OIZrqj9AqJa237rdbcACJlEFR6Yd4IhF6QmcxeuTfYomAp9WlhnCeXcZN6q
GgtXxQ6FsQvKjaS/gQVMF0P17JFWhnWWCp6vNcmSqAY3U6Z4THBXMUdNMTEp8WVC
ZvzqrQXYJrJ53nEx3ggOGM5vMVbYyvNCTCKD3bewzj6CBIQL1M/KxHk5xat7z01v
ghDauUPYTyU3zLQFL9SiXNHQpI/DPIMBs5ygeanpoJ84nJktZYeEIWVccBqvpS7o
6ba7zHvDnsNsJEMuPjWOkwzda3VBnnMGYROgK6sqVQwe+vSboPVxJVghuH0xhKyP
7WFUXhtJNLDbUDHUmM2aLAgajre1OpLCM2ZXh52IBhEArlxnE5iWaAnFDUGIAsMp
kHf7OKsaBBa1s/R932JNsvYKiClWHUeqTa++DQsE9BDmxSy0dvlAdXKs9tbRlSHj
ZGhbyfpgPLm5Xb+6hXz+HkaQGOX4ya/+timSAjBVjMy3LtASY0zrjzrgf7LEs/2L
FcKCvlrgP65FEsV9LflKPJOJV1QV1J3shFSJ8T3rZBOArRABCzVBcnZvZ8C9xw53
K6x74kpTrwaRLT+h32g4yJvbzazKx5g4rCmqCzfaUP3up38XFTRI+4pFs+nwSkG7
L/zOrMliWMVJs/m6wm5oaZP7l9H2KBLBOqqr0jC1fWYOPxOwPxBCO1H0khUXOYVr
t+v+wMCgJwd8qw97ipl3HlmpU/lKWtHQXkL6vP3SwHlmUDFyOiAQH3hukeaQx93K
P9I08hxbshsfAHo+TrGlXJ+IJChHOkahOHRF00rcQb9qqZXMzO8HsjCw/5GKuZZd
bmtvah68viWODLu5nBJVr+Lys+K5Ee8RBcjwp01F3en37wggB495I68HhCSaPzC2
1/uBSGW3A5J7U2oEkfIL25lyb+SlguTlbQdQA6xexxSjbIQNN8+hhM2cb27Pq1RA
HvEVoTLitph3MyHsHs5cpvbqRo1SCa7MjlUbbikoKv2ph0tk8d/CRScLPFpKoEei
EF57PQFJE/1e9eS1wsFwfxCGSnZEFd7QlVDby8FlAvSaiY1u1cXi2c3K50dtGcvF
K1iDrmXzOVzS6pdIN3Cky1so5ZH+a+ELjS8E/29Y9TVTfH+wcoJZ8uxYwOteS1u4
uNUz6mwEUJ89j2t83HSccNYoh/i9Me9+XEznBcc3sjdDO2/doh2bhe6DcnGOAmDE
hOCxHkLEK20hIjBpkGeJTwZC1DDgT0ERIk2FidoVavLzYPzYvoQOHW0z+xpAzFgv
RudzLFGchNv7F7zV28A3sWUy1OhizMKrvLttnU/BiZihwlHOsQbnUnn0E18SvFnP
ErNlGBKmRSbmpax3gDJbwiPADK0N415K/Jrq7LROIfqi3EVmvIJ1udpRWn6g4C46
oSiLw9nmEy2kQgHNzhL/xWAVD/IHy/3JI3oXu3eNswNrscLkdtUBqZXP8Xfyw+8Y
Uv+LBNPhFfhUzP0UJIsxrJSh/XtGGYxV7o3WOxYm/SAzsRvzQ4EMKD3A7rzonYjR
ZvEPGuODb4i/ysZibeeUqRHLb6pP7SroyzT1BMCfmTln0Jwa8SrWhc5Xgb8zWhLR
NDYMMFhgXcBcFeEicTWrVfwrAtI6KQUxSuDKH9dxLTJZ9aqxiM/fj0tV/xib51lH
iTk92NCf6qeY13/iy4yWqBYEeJw2T4/A7Q07nn87nHRPj0fI04mcVCnTP2gW/y9M
PtDbnPf6RQMxXiiV1lsJh1a//0pf9WQ1MKECJ03rfo+218K1EQnCT6B99TOk4lf/
T6OQzWqgB7s1UDvFXFI0k5FkiTT8NhlMK92ku2JoHdeJWO0xD/hx5ZGlcwapZPxi
ZfmBMm6e/7wStlh/PwYqOpgjLfsBwoK0QGtxD4gkUSmk7tXTBOZgn7IhLKMEiqkL
WH8Px+/TFA0zHZjcinxvhwu4tF4dhixs+TASL0bvtYNiGM/W5mg6Pm170mrSjHjx
7WovJeG2meOUhtGhn8wQx6BffFe9ZF3yL+R6m0+oAi7oIGfg8VpxX6nF4cJjj05K
XSmWRGKoRqts0ugTmBJcRIec2lmEmfpNjYukCdz/nNIZPFIErykMcO0iUr5UFpTs
1T67AYfF9qZli7gmbcnIz/tvDsTYtj8QtU+q9T7bgNjPd6Og74SSt82rOE7M8nWg
B0ZlNAvQa6pLV8dZqF+7wJAmKUn4Bs9g/g00XPjezqJKuj9F++UqVgKJ4hEU5maq
sfl6vV3xBd6OOHO2H/S1k90W/Zk2INH+r2reu0cBMEXSlFtrW2tKIDeV1T2kZSeL
RTJmbS9sH9v47wBiIkpsj+vTooILkQWyaXl8gPnqtLPuUhjN64/HcOfLC32wcgrx
rPGaewNdCSYCDO/7kOuDyhZbrxXXW4Xz8xUtK5+HWfm9YyWiwm6AfBMW/a9WDl8L
cWF0TBWeKj0LHWIBg9GEb4BDmQ2L/644Cv9Q5zk+5MOEY4nl0Jld0qjgUms+EjVh
IRSziCxbYtOxBsNQJyN8JsbtQZ87Rr86YulD2BmpAjcRbq0pz2WZHrcfkXa7Ocve
fa8NjQM9XctsidpSVHtSr3ZtiRVu9jLxRTS+C+VIDWkWqI4Zm+3nEQy1XzX6z6vX
EXeS+y8TAdTOewi1Qiv5yTMVS2h3V+RwsR5kwAAO9EZZ05cjrKLa1/eJ4BH6ixMf
ZTjvbh1o2mKA51A5OFa1nWO/Y+r7Kh/+XivdpzsALQkHh0PSu1fpSb1lx5iVtJUG
HOaiiopBiSp5/SVaJCRyyqS/7xbgZwnsHoorQ5giRnr3xMLXVLoZrogpYaD9+Pit
BiQ0AyWs/3wQOohhej1ix+bjs97sCi9iLCPlSvvGUJE5z06T+2g6b66vbAfIhTKG
KcIY8qASUgZQEVj6gITQ4AqNngY0I42m7SsMJ3iMkQQJ/LUbxwWU/fdfs8vqdbrp
IDRT4ctm4xv1LgsHuNkp/OB6Q/vtq5NDSk4PVJXwZUhqUaa+kbLXuqT/TKAOb5w7
fWxxyDtSqsQu9Y9TBNqUN2Dyo3/REwgYCXyobCWPBbR7fdyFFWROunM2MW8Y47AE
+kejPn1T/E8VT3suz7XKo4+tgNHZnhqKv8AvCordK+USA3zChTOGnmeb6vtm2gUY
Ig3SHhVLwugWd/YFWxsdujddbe7Dws8hm01/eddy00/PsVN19wPWUxZ3K66f5rG+
o6SLbIQCq6oqUQfvhvwchsJ2hnamXMSx1Sb/UzXMFyqxidSdJx8GU2dgdiCxwxPK
fxMDGcmjCOfiDT6xqN4zA1gtbno23byaG7iGBFaGL2nQHDBvCqgxGa/+AwbkBWna
c1oi+a9+85wOscRApmJGrgx339PlfOzmpOTAy8BekDtJiFc0Cp6UoCATgV9pDq1h
HMU8GGnuqL1L6LFvk9AD22zOrLHrZPnbcqxEU0JEbk2xb8jbj52AEMyf4oAhkUAu
7ZpRQ0Cxnwl86ardVuy57yI7Gv3tNm1sMiH6CyCvqJ14e0IQRzZX6ZXYCo3BG2bX
mweCXOsbivtTFvuQnynGrHwkLJRIFmA4Im9sa1t2bbAgxP4mO6e9d3CzkXB/4rgG
h5sTNJPZBjrGCmNjOxdF8OkPfJRAiW1/oTO7gKaeCAM5FdkKI6oEahj/x7yOl2/m
D+CoTsa5gxm424QCA6s9UQjJywmmrsqWmJJSRaWr9dj3V6d9DTWuqTh/IUe0HoWj
HkU3fsTPb+lHMndO3xMw0Kymtjp/+EGTh6Rbtbx+4ztqBq5TIZrC/IEEdC/fVDQd
7z0RQxUgECY19YxQ8xQS5AzeGsxim1ZW0i1wPpPLk9tQqNFYJSEKoObV5LEoM5F0
iduBoxl2JacnthZpT59zqBXpoEJyskolCO9DHKeZB5q9eTuuuicFR6gYqrJDwh5G
fUFhaYSlouJwH6Vdw+Igkpx2bGrHT+oxL9tWtV1N+H+T0jTzC1fcUjHvHbPPjJPS
hhTJdT4jXZdyrvMsmIzQmriFDRWw22RrWj1chX+ec6chg1m5OS7qxTJSnr3UbLIu
AK0P98tbvdPOM/hK5wJzkyj2GgxlduJUb5QQCnpw/TqRsK/u32rARele1vZPdRJR
A/IAJc4twTxmkQpoEA9f1X829VY1BtVqFfCQMKnblMXbnMZ0Lcqvcu+Rr7hKGeDi
xHLFJKgllwy+7j2vlIHJzhscCqIhiglYaJh6UTQRAS/d578wE+0bdtQA3KwOU9Xs
YEfC1+t5xQtH9fMZAlhB+cwvT2Qmmn7Rr+ttb19z+7iET8ybfZuJrWxQqovxj7Xk
j/IsBtyCrhJq0BEwjQXxPPD8leJmKSSDUIhlPudMA4O902Oqa++b1fVEhso5K6cZ
rA/nZwD04qNHIyEBib1ggnlb0SnhnRIaT+fRm9g/hJQIXNDVqTWe7OLguwAczcXJ
Lo7T+vdQ9eU4zpTUjgNJ5J0EdHJMYB4J+s//A7w8/oNtCMg0aANTo9piBuTLfSra
Uu/BG/F129u8pXTf4BaG0wq+f1DtjQT5I45Y0wSJTC3UmQ2BO04QB5nRpPb1T5d/
/0bFEB6PXHHF7XLrR+Uu63EOiI17MJG/9+4Mgizsx9i/LNU9gtMinHgRTWp8OwVk
eJ+Sow8ZIFFp/R2VdvdBiqMpI53z6KrAhWr9/Z28H3ztBLL0rBoKnuRc7LrhD5e/
9fBrInCwtCfFTb6teGMgBeYIHfW6b3K6kpYlKq6u12wUJJINESPfsjQWLxCoM45M
mOgoVpcfjKc2k8oRUlA4PHhr347vokRWlyAMk57vYEieS/uKMKwvj9cpvCUI/sT7
InGh+xOdLNG7LEUUKqYHzaqIzQXnUStazL8m+PKFkRcD8Zgfagt5Dq6iJutfQmiV
HO63ofDkgA5n0+P+neDgoF4651000Cg8dlTcjiE/lY4AZClK9M8lyjR+rXE/JNC9
U8edHCptuIhIS5RFh6pHtKyxPaRpyrUk2Q6BeJpTGc2U1kghc6DtaoGKuc5WT+WJ
jxcJ+n4A05APg2t45fJBV801kfzlWz7NuMZHH7TDwtpcblIJ+FdfBbYPKmR07BRF
VUJu03wjB7cDqb7PeFY8oW25KSilqRjwOpYRRqaLSWvY6vp9jA4soUCqRaw1AtQG
iaXIvWcyOCmrPMmlq8/hOktc7tIHC4ml4bY8UPck8vwK4twi30M89zTSXMfM/j0i
Giwdtkv7HBwchJ4X1dr2UwHOuHqtf+fpcTKKzqe+RDvThCdzdNbISWxUFBvezNTt
Zf/14QIQ1MnSKB1yZeQtstIgwdEaL3qFlc0tRwi0x6G66xqoRbA/kiueCfIS3IC8
P0wEeiFKXguQ4fomGc3Nwr+G91He15PPkpS5L8FOhSViGmGK2g4kYeKkBeJlFcwv
If1Fp3OWaPi2MNeRL3dleVQUU2tT6XnPrspftrDbMEl+mlpX6i1qHJap+LCLfzi0
MyQ42CiTMW13dMsQ/p2iFD9m1nqaP2UrpDdEj8gFyHr4zlvUuCaYWDAF7KI8YdVh
stGkHC/jEiKSpcsCXTFzmIClC/aEhCQW4n0I+hi/gAnaCgvRC+Di+pMJSoj2Rn25
EWrnuP4CFbVbFz9aJHkndAhW5SsIWlkSPRwsnZiBQMQXF4ME1V4H66wc7pd+YZ6S
D2kpjWPa7TrRy7tbixmbmR8zTjRdMHcX6Bal168nEfNzkUw25yM9BEdyxoWAEAV2
icKed8Is1dE+GIky7EaAFfrrntJv92qJUYVU/5uEZcwZXx04BpjNCi34KoX1qfIA
dahLMBPNfB0nI7TE/m4yohT5yXTzKHWdN98dN5odZ3sTFFox9GjW6QGuxgcpYBnX
AY7/GBNeKRI30tU01rMrUoLDKNO5fcPUcifohWwqyaBgFumVG0+X2dgSSmage/Ob
NVeRpOhbFnN8Ygg6rGGk2iBkK/swUXog7WNhR+7d5yUT/a4uxXQR6eP0LxPHZzQ0
MmmdkXO1MOXnoakNXYsWlajICfrRtgSF2LmMwA5uKX/7VvMFmbsnBcbFyZlKZfr0
7mZwIhtDEno/1v8dtT2bT/CQCUYPDTHQR3UQG+MTRSzdvgyfUokmj1y2t9vPS9l0
2T3ZKK9Y8RqjGxMMjzh6gdBO4tngNne0bqGYfrCzWL3/IoS6RWXJwDbXuJqJf9xe
JPd5gmJDRwyUBqRxSQ9ev/9URLSvYqmwzVtI015R5UrbZzVNgBKQfxevVdaYtvdl
SXkhT+ihWTJpIxybBHMEe01/cRZsnFrohA+BdzXwG3vVtATCpIioMV99bu6rlbro
NvsDUwcuZqdnPtGVAf+dxwUqfMUKTKQ0V10vzzWIAJ9itlDhXhyUUsmuOmT6RXXX
XlIWSaSx0iwyxy9pLlbgL/wnJOjv+hW9MMd3886usZJwT+bnMDaBL2lGB3V2PX+Y
QHT6mkb0Je6RLyOXAhjK7jfFMxyjAPvGcR5ifEdMvVXMt2YpviTL2revodwWh7FY
in9RtxHgaU0++91LdrnOG48WYbuG7tFhpurEzbvra1eKDZ4ouEgPmR+3ETiP37c2
cI51uWVt0uwpbU2HfhPVzaz+zP5XoMlYCqf0q3Uk+UL2rJkLdCGaS+rlBL1LevjP
miROLo4hrQkRu8jpcfN3ksx7uIOj6Rt9sLQq9fyE1UqE+7wpJEtdGbv1fcyf95Xf
WJaQ9+3tZOckkkOS8I6F6NzLY+yIHERHLc2HwYfWm2QAi7CCCdc2xpIl3fRKej2O
3QKyzOJM7UTCDPwZyK8JBbSzdkTzWeHU/udwkM0gwsSqBNhombWhAQ9++oFhzw5L
Lo0gUK0AV+W5tA9FnGaDpb5q2U2b2wLXEdOP9qrYuI/Fpni+snml2HrFcjlDVSZ2
PhRPP7GOVAAnPS87G3yHANWsI2v7FJ7HRP/bHHhszJQuQT5d9VwAJBI0bvTxNrCW
Ea1lD1LRq+NGEpKZDynH1zyN6DoYbQR/LoaAUPa2DkY//uj5mD6ObdGlb+v29Uep
6zkqAj8BlVGbMY2SxdgzaKUopR+yInpOgFJhBU24uDSY84tHfpilXPvhPT0Gg1oQ
asiGkRRzhPHSTQ+8YZj0EoAC0HdXP7u5L4+oiGdYu++Z0B7WwGoyi/tWDYyU188J
6zHPyN7lyFdlTHGTvVFrPzBp1KTNpuIn/sL+/uvnHkY5D8LulbeW8P9IiNmQ/aO5
dswRpRUimOyTU3mfBOVpdwjb1c5XDeh3jVIKNv8iQNOzTTVABeAG3qdF5PEI8gzL
m6BJaQbBZgKh6AfcnxJVs7zL9qkmVhAP18kTIK/qz/ryMKJm2TP3IlBF26uI43QD
3QwTN10hnCpoVMMBcn6SJWNNFNZkZuxXk3UHAOqNS2Tk4zZNtrznggfsohtXlLgS
ZN63zg7Vda7kGTj4wJP8Vvug1rzdlpgnJoDAybtU3LzgEUjgrKEmheYS4I1RmiKH
QJYPo4IyN/2TZR2QrQwkaYLZlgaEWp994v7hYw4aTp5gWa2a5aHabpIgFlEXdWE1
bNbX3wsmX5N2FTQ57gCOypFxtotPNNd2ayrdQSBbyk64myNl/b0ud/QQ+D1SyCZM
qoW0/YZM8K69s2NCTuctIelK9MRj79UjlKqNPp3/p1c+KC/q0+SWKVzBmaBuEXhg
Noto1gp3zhen+Hc8VpT6mHR/GmV9/2TAxONdrQEHDfSdScID2PPBpsOEIJtOaKY6
1WZPTQo5/q72HWo7qxES4SthAN1FRR0gKYfA3St4TDNEULlmH5FBNEw2MDzajVUy
yQJf2xKSR5f3z4haNw1bAXGMGokyOYafsoLiV8IRUSwHjESGLZNgSh6IUF5uFPd2
xO4yQnNV/0ndp7kS+gUy3yEQJeLapJHz+MYPl4rJ2eNZWagOHcomMMqTuyjlbsnx
RWQ7huth+N7YOQDOSGXynvGIRQX+vBKwBTRIzyjnizIfcy6gWDZqYNllU4SiPxdd
O4ByFJrW3ntbvpSp73dkdc1wneattwBpbIxHETmiI0pCI61a1vWE/KThsm8HomYi
/UiaU8omtysGdFRUmXXAIUp23SZqbKoCmDxb3pEI0SrQz2t0KYJVi6ZkG7K9O0V7
azF22RSvWX+BLJn5enZDspz4TW+9vRpfU9GIs/F4+S+gIv80WC3GHHs33YQX6Nsg
kBWBdkl4HzjMptQXl01vEHVoSktiuHkPG6Z7H+XZovmq42GNNRyaT5m1zirCutSo
NXG1+Dq8+fmRNVHRPkJlCaS3LoMFw8UVX+UO/QXY8HJ/yvqs9S1SCy4VCI/F9SMl
quNQVbHGHD3rtFrdmMa6uM6BquZHJN8P4VFzviPZ1TVw0AkJ1g4BpkdZ3DGT0g62
MYnkymlO1IgHWVEy5N9UIoDmGeXHfxqt0RGwDRHyhDhe/66mRdeZqRhRFLCZ8FI2
DQNkTR1MN/E6MOHNXTJq6bI1zDRJPd0Woo/y/Tv9XzsrF5MRDu52LZnuAfRYykXX
ChsmDXFxZEPUlNWjTExzI5liNZPkRweEo6wh3lle1HbRrqLUK2o0JN1mvbFhaMd/
bOjzEkEjckflAJ8ycBI30PTQVAK8FYroSvRF+jX5kka9tDoPgovCBZNfyN5ovsuH
LISB3LzAi4ICf8JSi/+jzuTwVQtf9TtzUGm2ERDE3vNUyc/sgV6haK1UqeteCT0F
GKnxrxZB2IFyp+gSH6PYSK+ZcJXoELdm2RqzCc5/59js0aNt54Cc+7vfgQuWdcPg
YxUc9j9oICVn5yHCD0M0+HwKTqAlexkntgYNkyuRhBl9nAlZkxQUWWwGpoN7OkIL
c3yB6t5p0gDioNER6gElP/3YqRbKyqB1Q84mER+htECUARkzjtQyqV7yGXZHA1ND
ElYhpeWFI57MKvmEsPbUuuJYtMk0rRQUg2+IeaZiJalPc8S583qCNFhrrQt6kFud
1SpNOPWUMwdhX5F5OP0reOyZMdFq1WIisIzhWfNtlF3ZEVlD8FB4ATHBBmerUldJ
E69a/J2FIAT5pNEOtUmDsdhDoHQ8cvD2B2CGALFKRoUehhCoIpAz8wybTkoT4iHG
S3SocYudRqUEs+6Z7ToWU+Y/zLdPF1zBUFqDz2OWim5EYDa7Qk0DQfXYUYI53dkQ
qD4TmYR/jlKB4iFgIDTiGqnCMjExXB4IpAuiAVI8F06ivbpTLgMKSDsN76yaHceU
l1xToNwXe2AzI/iGo3VtE11QjC2iFC1UUQzO29LBdqtpOAZFuqJJzEZc36ST0pNM
fTWshF/33+IZXFu6FW4kd9Bui1vOtnLiKyxxUv6YfJSDXDqu0NovNpTfPaxmzbd4
hSoX56U6U7O/GjUakrrJZKhTjP3pKg1hiWPUdnVKJPHdG3226KGIJNZdzLwmhwsg
UDItqrrhzPN6/zys6niqKaOg18z1IRovwkztlNRWncSBoCODRcfHbnVBdeFoWFVH
zBoj8advanw7wBPvu9YfIVRUnrLut9x+rifpsHHl7NZEMWjLS5hVCrZ5Z+HpHu25
amgAIAC0FKEFfqgVqU+jzowdRl/ozuSIYjTRj+cFAgB4JcGbZbRSRG2vmJfFjK0j
aCOS6ooSVsoquZKLAVXyMMYVjLoROiZniTuPsqvNNe8KJsklY4GUDhqv632bVMg2
W0ljnJ+3MlgBiIRZyS2YAZiUPb4ZqjVWk28P3EMAvEP2Wlez6vApPxp8WO11VZLo
Wh2N0Ro27wRbCtNMdj4OZjABcqUZcIk8wCF1JX7+Iau2YDXSSDfcledlPdXvbT/h
XoLCf/OwExVmakuVXAjw1NJmCwK4KFBET0HNGLTLeUKN/NRn3YGgHY8gEFgfmbf/
ROc8AcgYNpoBXZHOxzWjXJdvrmyDCc2P3x44MdJm0aSv7pq95DtnvOhKoHwOqAXA
B2LmodrpwHqbfXuKrR5DhoiZeudIWXGNZXOEXa4wztUITr5sH/bxtGtjV716EUiy
jadBOPlnHehaP1Y8CflBa9zYWFYHG0zw5/XyQEo8ps0eH5dZYyaZjRHt+ty6UeFM
Lc53fC5Xllvbm7AfeTdqRhY7tj58rDMgDQmlxa2YIhFzMB5jzky0JuREqmpYJD4U
VVL0timYF9ZS3+jXxGOp9Fim4UtpLbZfJzTKXsdy8nKIlxxzUtV5OZfPkCn113nC
cbxPIL4Fzzn8kT4SnlfHej4NmyFN9yVVEXVAnCdSn+TknE/Ou5t555Z0os42K/PR
2IEoTOsJ9dh/prNY+jc0QUgSFZDdsFhF5D4NKrHPwklVKCLWN3lyaJu25XcnUkOp
2P8B1zJyexpjXjBJ8MUu1b16I4gnS6yI4pwDBYxj8ln9cokBfN8cpjtTSSivUPaF
S2H0sZPL4D4TmTjo+oofWHBAnwXVJyHbwLb5fA9dcMeH8xFuXbRrjLu/SS27fpkm
4qwnqqSipYarxwifKk82JcAUV/e8Xwf783eboIh+Fg88M3xdmk1bNmjVUKxaAFHF
tsKzgYcQWgtJLPV6tk4TI5eGVFWYVPnGml0bjE7Cx5p+B4NSCEYVoCzhDMKZl68I
U0Hau0n3bEivX5n03QqtQi7L6E4aAoEE91Sh51TtjlfALelm24bmVTK6C9k9l+i7
AIJjRQzmAW77mjhSkN6sLXP0X9GN2vhOw4l2XAh4ZTFnlEHbQD9HlG4gy3i9rr/p
inoqzkc32IT1WFUjfbgSKYRxSNyob4Ep6moJwgZsme/uj2yRyl21C/e6n8bbvnd3
Ruz45j0M/z6Vva8a+YamCTkR8q86FeSqkjS7CzMqaFIGQbN3ALZfYBNQ0/22ss6o
tnRSNe/lUwFgOS1MSy4lFc7bKar2DsgP/thbwhyDaOOJUzFR4eGqzQmhcTWY8uiC
rgki1hLgLi2kQPyeusBydZmEr7PBFTveK2HoKc5srHBQNbIaBwp2cSdxNtYACggI
YqX7eqy8/aaOPK9RShdDta/06DZmlh+e3eKwEApyKwmPYDMSj31XwaeZdwqbcgrn
3TOVDXIa5Y8taBUFM4ygH/25FyXsd4yXJhD15B/AsCPjaCXQE2lIFatv7ie4sW2T
9BTioZ+YxuH2IDz5iSCfPoKSYK6N/w+m2eFGobxvltle+KfSufYNm7CVrF2pwmWc
ZtmPeeFaKTUCNFGkgM15logO0ObHVEH+VgSSpPTaOS4gHFkyYTOJI/RMh16Etdtq
/yVEsUhjLe66jefPRjICAQZvaEMzsYQd5ad7YXugWqWreMVfaj4jrz5A2CsGmL6g
CYmydaq+W+iVSOjQXxavsSl9DsSoJYtclCvTNtL8qxPe/Orepm9SZgvOVdvjtkeF
r858daSgbkmTG8cAEd3OvHeTV+T1q5923vivMRc579wkyTgwNisGyz0A16wv+qvS
KWWV9NDfYjZwFhrJ+bE5ILeKugBHBguddfkSvUw9AD1DYATh3voY1+YCJJ1NmgYk
BR3jckv0XehW2kVvbTi2fkdHrMqxHdkqzZZYFC63avly0w9YzCjwQvCLxhP1pFcG
qg0RzYQ/6GekVWybUFhP5I5nERBRVQVTaYyr3EmRaU4SJkZh7jZsN5Odp5pjaGSY
/HuF/puqFW70yaqae8sxA/8afOOFDRqXag67zkM4fB0NxZi9bCNIDCsnRRDRAquc
7WnxF35jOr58B9B9NrKmSnCKgdr0V7WXLLQZH+SuhfQx6S3yM94PvRZBphRT9e3X
AUkya00WLvTIqnUrJF6rvLHgpEzpR9KVH1pFu23layKn4fldZQEQEd3MWVa3MSUD
SBlJ5sYOuC86ZCzFOGX2ZKs+gjAuilh6yyS29WHUplfIvKgH8kMIv8CntAxsHqg1
Ok+akm8+geTD927RfoiaVAzPiiCG2FcoJBgLRjER5Lqj7jFa4R3mz0ACt2hW680+
8NW87hyo9sc0CbLVUHrbPjOWeydye2t6Ghzo2abMLb2IaC7QQICspyd0YxFNIo8Z
gSRcZKUQV+GrjVi1E6rzodjlHD739EQHBlfauko2Y0aJbC4+FndyqFP1glANR5Ba
RaeGQciTnLFV5hWbyVr3gzOu1SAEqwtCdF4fM9Wlzr4Z2dJEGxlh0iGuvLzikpH9
7rjwbmfSsHRlUb4Vqm//inuKutD/wgpIl6vNIx6KNHEM3+83nuEyXA2IoTGzuXRX
a8gyC7W3d5sS5PD2+ZcuzesHqGp2NzJl5QobtbfN01q+lQdqHByLfa+WEA/mkhal
VKzoVx5lrwO3gyacUVsrdutDJWL0nUuB54Axgih0cKIStIjy3fuzTXXItX8YEg88
hgrE9fOlHHfsnwH+HxMUfc060PpiAh+WfajPKijHqOGboj9CTQrMZaPACjfZlz2C
ub3fwQ0TxmRzcHfdb8eXsyBzrD+E2t7IEcv/tHsAlQ0aOwbhCCLbj0nG8VzIAoda
7WWZE/Db3gaHuPDNhHrY7gr7Cp1j3q7sQpEC+QJkU73950p3zscPsFRtdprVc5BI
UYlHG653/7SP/enD9Ly8sInwz/Ry+caQY1vP06v3mJA2dmMVWvDQN6koHw+Jtuz0
g3hQiOHR6aErurXa9nfdWnmP0dzEAqzTE70pIW8eejeaoRKE69f/SCu+6Xgb6G4H
Io/uZahAiSyAf0csKXRVkPUyYvPVNFGoEvxPF+TlzzJhqAmsAkpTQjnv6hwxaAme
DFSqjnd5LwD8eDskS+ILz259P79Wq8soZ5OHkcl0RT7ict5ge5Oj/AevN3o1FdBP
7FwF28PV+pSiORRk9LZxThKMA/9a/AEmA3N0gMcSs6lxX5N0kFqnZxUD6bC043/k
SXL5jG76D9aUtSvLmxbrZtx1/VRbeMgRSTBL3ZNsQgLnkXEDgxBKsQ7xByzvz4s6
Md2cjRsGSF8C9R+/FMU5ZAKFTNjl/tNB9QaDs3NXCLe4JURqBHjo7/zhgmUe92/v
xcFLa45+EyxCdi+sUeliOxWwWOfDz9XyjZVDk1nK9Mx3hdbDXti41um7rX9hfWrY
VQga/zrnLsomrdw5sGtMiq9+HNbG5Jc8EHSJKa1T8M+4E8gn/KHakY67q/iV7Nc+
633ShhC0ySo8qf9aT/638OyxCb5qRBko/omE4+lm5BPpowR4lgAJ0rBbrMuIJkTX
DKDFZXOJk8wl/W0tojPDos2vfYH3VD1pRK5i4zz/miHUZtBujcixTvaRGLZkj2ff
kKdGgTwQfz+TGhsV9ihmqk1bstHFIilxEd9L+4oZXaf4P/V5IwUUB2ix+do3key+
wOL76T+EwAgiZCcTjbmjmcnhmmRRnrsuEEa6EFWl4m8tWfAif75SP76sDjkxhlo3
McoU/XX9URf6PBxxPRCSENzle46tfrbznpoB6FrHTfki9rBdJ8LnpaS2yafRw/B3
cMhZrOb1rik9TMvwRJUwuMRKMWCcP7Guv8CLzCoM4MS92CeTe7Qj25pE3Xb/GMHc
UXO9O43zYHUh530fQXHcsXh3K6J19COa4qzVdIICxiJNegAN9wFSBWg53NMPZ6nU
RGCjMs48mWCl9K4PaAXo3rcA04NP1q/wKEq6hLEBGixFh7A1w30ukSxdYDSv4FLT
HKX3b46nNZh3QJyofaDIE8HcQFwEzkDkNsbXqfPW50A1aKyDVYy0a5/p8BZ7MAn8
zW2cLFq5PTr5SYKq1rDui4/azlOlPnW8N7egyJfYdxpdScvSM2X036LquvVl8aoc
KS5km35VRB7PPJQeH9LO6v58g1MFM+qUtJN31rncxDaIoVEer7Kxr5YVdLF8OZpY
Sv/BokYfsMsfRJAx8VS0Hqq2A8aFOZG9AZfX1qctZmeKb0Qn5d72f+1h6t4jXfcc
dApTAq5AKiGWMJ3aR2macMaGlCM/gMFv/gyAFxYnrv32DqpO7oLKXnMjHSsA/XYO
OPj1BlJaTO12rHgq6crgL00yZnczmBoV1WaT2++iwSrfFobhym6Hi9EK1TtBhmY7
VtSYe4e0R9v3gU0VVNGIP7u9VN1RLpCS5MPl++RSonBD3JFcoMbxqe9d4we6CnZc
/32HDAdJgS/l8i1MY0s/sqr+4SVM6dnMYWaaIbuG3N2cra00qdFg05I7Yu/zZC0L
qc56tyBGZxflUOm1R9A/J3REQ55aJt6NMo2uIqX2o2xcFSA5icqUmcssnmtum7Mo
I7NMDUze/LtFdTlC452NdXI6os6s4l/PjgHY7/fZCeQjOqLB1jpr1ZZxpdMHo7gn
62iczWyXJd6zNltWvOcFWjvmZILL3SpO8/CcTkdKTpGjCxRsA3d+S8yf8qGyAbCE
lKFd01k46sA8uvVtYOrq0d7LZT5QfdCSxAcow2YnOcVFcSkq64uFzHFddY2AM9tm
5wB/Clr7ZhkGVYVZXdAqYVHE0afH5FQmxq+K9npOAVSJyRmENmueIhJrBgfkEued
s+VFNA/t0di0GSolR9EDaQrnW2bVZ5qDt18XALLUyrpEjYMzJ9togOgKLaaQEjyB
DVAc8tdCYLtbvNzcm0UPUrlZ+ERb+wWtROgEh6IbD4i8LOXKvukTBwvaFYonlY9G
1bk7Mx/WwZU2oTpsBZYYAgPiH1hOjeCdBGfh/VhMAvaXUi4y3/TMCsg0XjDc/3wy
ikpWxiffytZkqvfLqaqjoxuBi4hmVauPlX6tf+ifLhFjzvIUAhXEB4t3/lo9hUiY
if8U3GzcX35hHwNTJ3x5RdKvoPy5vh9svmhD5uOzjv1nsOaj4MIIVLP9he6iP1wA
U6/joKWcK2QD4VVk6aV9wU+D2bzVcxj9p5mXiCK59PrLXbbniDqIcpyXFYBDTkdO
RgfikSqba70jxee+US4t7d5wLs4pd8xX0Q9ZKR/uLbtGdnAoMeKR6Ej4bXVWmPM5
8QTLuBwYGDQ7i1pjZu24M9zgCQK1nFDEvyWOlcpJcStmDYHPEGepf+++M6PbnE5U
El+Htj4wG3wOwt9jQTQbUEszUivNmXH/8Oq5EfQNQilv+fP0qXywRkER5vDIzkMv
K2O3zMvrWrU/yxxJIKXJ/iI+JcRI17FhLATzfJF3hIPxNgca7Jt1FVkpno4mVKQq
IO6VqB4BhJBmN5TueaJx9eOjDdmXr3Te1nsmqNmYywd1jAbFZ9tUq+QGNzgWhVO8
HWzBv8gcGmRZwJsSUErW39ohIH8FA6xOBnWB7UwFQ58uGtHB/SNCZWqci87rDCAn
D4wJmJC54udI+PYL3+wYlMekg6ZWLKhFcDBKIr7HednTs/7EaqzlOupn7eV2YeQ7
m41nXkTU6potyXbC6Av3lCwgyonIjsqYv8k9qEIXqtMD5kg1Pr2z3/9DuzLH5TGt
vAQAcuxVIHT1km8N/pow2srmKKzH5oZkf4OwHA0Mq+8P+ekcgJKFsijaywIpIiUg
8xt1mAbDwfmfV5KuQ+Y7D9mtfjWd7y0ZdbSpm0jr52eZN0dQ0XpWKOCG6yd4RgQ7
lQ8w/aYM9Jgd2kjKfJUfzi57gRwJypsYd7MJEyct2NDEdo/Sr8Eevt1qkPB1X+tO
0TAd6ZtucCda/ryWjGNGKtLjGTLaGrZtp59Ur3i3wJcKn25JzQHEsZSQ2nY3Zv/o
Uor++jFGc34NLHogFED9Rx5l4QopZkLNdb6Zo9ObNpWTXiipeu6ZpEFnEojA7/XS
WfJx8yf+ZIHE2w/DbvkzArOdifmL8FPzpcECQBZcwvM5YVbDkTqnTPSFKG/yt7Ev
bUg0hgG+vzkW2tqCAfvvOkIm+QjbYtmD5drEGmE1T8V2jAAvfSx5SinXqTINfb61
RxEX+mUTGll5//5B5lmbrPCuG24fxtV+qioD02a3UP8p0fdsdSI6MHrVqz+fBY+B
rpDNW6aTzb+QW2S4dAp4ne4jtma4p8IbBesH065ePpdxxHZPtdm1iZRpla2sm0Ta
62VtZWBeXMFlNlNCTdcsNcHhRHHAIdGQqTkkaFTAhFLXs4PvXE6NXydRjHu0G2YR
Xm+L3Jgi48rwnP3QaPESYtGHN+fMd7oq3RbwsYC1tupHA/VlFTmb9+ft3SMpD031
j9vGvBOYe5z9qkYBH3hYX/CfyOQDoYe11w8IIsGDxhn4Zggn/K8C54gQoDct+AWZ
fViwJbUI3qzG6HvuKPoVSVVSkNuADxx/bOxQflnFJ5NZihcEyohITiFvRgjq4ZH5
T8/Yfe8Cox5YSD4c6ZAKJe4IzM4b3rmGnHRWjo3xvlUroS8d2E6y73Myudz+24PO
MJXVJaGivezsu0Blc6Ipo51CvYyT/uKL7mPweq7S+ocW/RmDQBHXqGOcuoeMgmgz
EGPnvK6AEwkGse/j2k8JVjyJp0W01R8D/K9QTHhyqztyNYsYEe67YeXKUZP9XgH9
eu6dP8/bdhKI6m7Aq6NXwKSt22Ar912LZZ0tGxcq6TpbJfceN5HZARdyxBY294uq
pZexdj/gjnMUebfBpIOJukn5SrH8j27ZtivNz06bzzeU2CPZew9Evh5dVmzd7upD
4f8gyuro8sj27VdnX2XMW6c7DR0sT8lb3wWsp+b5tGvjHr6tjn5BzBif9vcb1wSq
pk/kokG+uPiJoGw2WJ96SJgrGY2UYS02RSYtKVtlnZkCvACWtRmofr/d/HA6wNws
d4WWUjh+CaKz5Ehu6ovMTD9wVf7aMXCsehMr0jtoEisEjOpnDQYKSy+QKRzZ3dDb
ibbYRKMMzJNK+uEIw8hNZ9aFSzRLxfQUncPMMj5+CqT2058me6OwEmtVQ7vryIix
/CW71Vs+YePIvcUko2gtR4vYEpraivaZx67StbamYZgBQkbyucpGJiNBNKfPNmLz
KaIIi54gZiWiG/kPbzzOawdxUbC/PVfSOCBjarMXSOhbUGZMl1Bj2EAEBicfEKAE
wvjIS28lA0cfbAJhdOMao/3lrKG4Nrcc6iHPghPqCwVcw3PVTTbXlChRyV+pvins
U0b7xhgLTrTGfj8tHsZnEBi9RkIBtwgZJG5JRhjcoHOliBpqFjX3zqCsx59YG+sf
z01RRc4UT5zc54k9goS27CjEweA3RACF/Q60qd98MTU1BJ0m0BbWfx66D/k0JlJf
dTtLN5jza86ghSuf7KtGIrvzs7GXHOnZqGR9yY9cJJdXQ8Rm1ff+OmP84LytS0uF
UUEMi2OBv1yD4p56JXoqIvszp6NQ+6mSEtQmyV+3tu9um4CoBImDqOElnJs6rWzm
PUF6RqkPYjicwA94NIv7QwioDWLHwv3xkV0MPcDZ/zDNmwXJSAG2N1ozf6I8UbwR
34TJlizUGBrt2vNNxDUhVmmfo1xexUdNJK/nYYuKOVL+6Vn5/UosVjkMj/RNmche
sl9eW3cI3E/arjEoUyb2dU/X1rcyXR5k2nIWTjlwZF9UaYq2GsWaprTxzQD8oJeU
aL5RiOoSEaBVjYIIn8WIL07Pgka6q21dOvKu2/CWno3knOl60UWbaZS6je312cB8
aSW6i8JVwz90Oc6h5LD/GnncdM8YBVMe+20UWOEZ2cJXtiCPDXR7P7xH0dsDZTLs
M0NkEBRk6eek2zV6zLX0jcgncpYkwFsjsA2r1IkWsIfRha06rrvVXYZdDYBqTJef
eWWVeoA8avdsZh/MnTi39dwoRZYRgsuIusgc//YRd/SKEb4tRF4wrTGjwCt9zLFy
mRLneKV6+hpIVmkuaexjW3JrYPV9HtNnTuyZbf/trolLWLZxoVpDa/lDwwpiFRZm
rgS5gxW+lPmL/CviltL1/zjIj2HMsdMU/SrQ9HfXWSDwxRK9JjosnjCD0Z8jIaD0
ugou3MPUcNvkdomt7pq64SOcEaDDTMzyv9mgFFMpgQno2ZsmogMMgojZ7xIBW0UE
/Wv1eXcihFGpIzuW9j6/C5LUMwsBxGQzXAiVbyEXgb4pEqI1WZi6OE5fKnlyr/lj
wUQ6t/PlAMjMraAL8jok4x6QD1cRVsad1NcQRuWnia8rX612iCyRGWQUip3cDxSp
okGtzdr6vMpIS+6PBjX23bK6q6wtw90G1Z7DqUhNk/VcX9oQ6Q5FjEkN4jOWtlci
f0A9TjD5GF9G0GkvMT36HY5TgtmW3L4IUhDcGGPAIkTqSQvVz3xfe6UU/hRQ94Wk
oTRTqJjc+yNE+DCsaliwa3filEykPeif2OSPRTxVHt9GMNRtTI/Aa7/Sswf1w1fF
GHd2Uo/tQ384OmzF/rqT94RJDAOTJu/VT1dpcRH++IUBP8fGF4ntFEONgqDuXVsn
xMCX3UzsHTEK5EGv/hyxctyT8h1yXGFiuNhQ8c3Xn3zMC9IilkFq+G0NQ45ZNgV5
O45zVHHRXyItqLUxMfaM386k+59ANW5fbumHhbLi4EaA0QwQ3g7k6AyWwfg4K4D6
xZ1jFuZ85l12yulh/a2Z2SOCG0p7wuuYXviXe6rGLgQ7iNslfVD7YkDTl4D8ic0w
42oMlDm5VHUx2HTe3Mgeljzk7F+KDg9MDrilLvU9HVts4co2GQCs6Gzy3RTpYAdC
7mBJcYiex24c0oRX9JNZvPxsLQWkPRk4/sUpk0pHd8nwEmt4DKMM9JUr4RfSl2rr
hZ9yPl6xUJ3B7bvWKcRik19oXKXkMncaaIDhOjEFccMiWBgf47mEUjIXS0QS68C3
1ZQYzQcR31gfHs4Y7LpkUQGKaR9ZDN8tkfX8vWjVrjBLHfJ3vkNbblvj3Up08qiM
iT0QNiXVXSFnUmTsqT59kzknP267fXV0K6Tr4q3ONhMefWNHIgD+L78Eg8NyDAsY
lKE2WRO+yCHqN1N0Qes74eIvPtQigaDY7t3Evqq5BRFDuobNQVDazeRpXJg1Wjjd
WeqY1ainvZ25ymaCpFBTqjEqUw4vNmSNO2UpcL1IfVFkC+pQ5iEp3w8bHOWO0/i4
GqNjpK6n7nW/US3vzMWTKx7zf/L9RONnrqiStcCI/jJP7bJejYwKXAWaI2AcuLZ9
EuNoZLZpZpxyg9zroqnmd4a6c5QGKQv0FNMVRlzvdu0MkfNOdX5SDg0PHOSVD+v6
IZdaPAwCjRwoCfaT8Ndk9b8IpiCZaBxiNaUtpZWJvpRxoujol14MzVMerigZW8h0
Kk3cRLVBJOIPUfmN4ti84cRDUptjOkTsl7sDh/H+97jNO/efpxdQMlnU92udzd5V
BvG4/wTjc1gYNzEOvn/73lL5aOGTLmVRgmgiMjMGaPfklQ1dXvW7X3ixSJVaToj0
7BzCJ7ubpcXAiGVNNoVpHQwdaJwbHtW1oOLUSxhWp79P8eD6G273LPHe4tjziNEA
nNopBgjEV9KuvF7NeS/46TcpDIkbnJ3ka/aVEVpUtS+E2XnnGrZ6AmPiF68YqHGo
oLhWQDeaMAgSxhZ279bgb2n/bViQhp6qGEm7Yq1twy8eZ9YZqCH6rjBIjaofAcDM
cFA+LJFFcFYN1lSne2Bw0YYFu/ep2dTJ30htjltaYIT1m8pe/jMANst6Uxo0ipAo
gLfnHIWNHVljxeEY2PKJ1Zn9+Vwui+GB/UvcLblVPgWYJeaseda22IgoC/qupmHt
nivNIUxipCNWBBTIQuKCftIopJaQlbq/I9mFJsJv4EstqzxJmcN7X1bhRIEMbfRv
xH+PIgmrCOLlVN6IDWxl2wBR1sr5ibOL9pEWqDhUGMY44VGtQOe69n1etx3b4rdV
RwhM+nosas56xPWb3nY2hEwzMymS5L/He9Mwih25cNftsWBgVUX6Ky+DkPTr5iPN
vuLF2+Gk3vSxm7LMfsBQDWf5ZK9JL4jRcR1Rpq1X+8PrAmrzbOZmrYTyguNLfXmw
YMWz5CnkMX+gNV9MeEtFUDU1/al75NoesmJQDl2CRTBDDHSL2O7mJwqfx6HU6EIE
T8xO4uz/NT0/1mWpSEDRFsjXIe4VpII0bhKwAPPgNOG1M7dYWGueOTq8Kh85Usf9
ixxi9yI6wrIuarW8AYM2HF2O7IfJVtnv241Pbh5V3MpMCGm6+MD31h0fkBBUMbyY
bRRLUzse+DD53V1MqSW6ERuOsP0za7FcYbRbPK9xVw6eJheOGCD5xXBuM2K2XfN4
QLjgzFvgainvzZ3Cb4wd0O0XYkawXztWrGQpradagOKGo7AHDSr6rTZ9p3RSRfWM
A2SSKrSSxs5LeCrDScGfRYdwJoN/m8wA9olbu/xvojFe32VukdZyLekP91CW6Ipq
Eb22980bq9rI1cMWhF9+X/CWuVhJg+h2L3L4RfT0LABjmLQyk4lPgHUqvCa80keJ
Fm9WU0qbp74tudaSTSlls84QDpesFJmbh8wTPcpq1eSHgX6QDWsD5S3TEPcsZecv
DuWb78S7JrTZwD2374HAAWWKSBkA5gjZuZsg8dVmyvjP7PeeuUhCQ6QgfR/V6VNE
+i2vY2S0l15/vre8fmgoAaQuqQ6AgN2mw+jBb3/0GEGLF4lO2zHOmNrRhfx+nnBT
hh7K9CulJxWZnnxGumxrYRDyQJACRRaW4SGPk0YNFUlGFcwiWmgxnUCRZdrkkto0
g08yjXLvpRPjTsLEy0RV1SPfi0bGh4mEM36CFCyeW19y9k3Q0d9DzAWGkZ6km+Tt
9yFLbV21DqRCIT3XNiReaYJCt0rE+mn3TqiZat236OwAg7REQ6F9TuDrH8Hx8sf1
UtO94/e9/XdwCQj/sKqcGN1dyYoDjpKrzvA8jjSZyv0xIUWZN8k1TPYxWwoJtvDB
3/vurj33s0D98b9YQycynLIdAiQmUe4pfXhP/JOiGhlIdHbksxW7yFcNFS7nyHXk
PVfZ/gQy9ipR+/D9aB4LHQarbsYsOLXV1GJw39hD+hDDV6NDML8K+fiTaU6O8BwK
xhzb95Z0neqnFcuixIdIOfI0/cS0eFehxAEOLgY84CKgcVJB0QTIxi5YhHE83vuq
Dcewv3/6BTkI3sOYuLWHqsqG+Ln6+rLP0NcjQxzGkLhsqT9Tc25C4b0hpe7TqDT5
7TuI1eP+hImxhy5J/tSQsYJX9VOJ0aDERvJVqeMp+T8acA9pce7W24/3ZhLIuuJW
DBwlliziSZk6u46flY50OAvr5sYIad1Z428yI1RTSU4HqMRLSMDwbyBG/jMPLXFY
U3XQ31dXzFKDHPRDNKiAtmzMt/UgBvAT5IUFkiHz/PheViAo4OpOqLK2PEx7VDs9
oA5XrSEsrWBoYRRAaCIXn3TquHKREF4I0qNHeqa1GUSe5hPiwY9bgrP7UWMUZ28W
UcsSMaD5IiRT0k8bEoc6mw8NUGMAEr87ynRoePQ7dh2mwdF0EahZXNlLzn2o3P80
ZbI3aTDRrbYlIGF48vGrIbeld4HoUUudISqK1ckGLONN0hVVGUFkKe6D6HM0//Cn
pXCyb78xaNMQ6swMy6TzHClJfnSxabXABNlwjcwPRKVT4KTP9rUxw7zhJIEj5x6/
x//NztS7A6Nqil4HiU4YQ3sYiaLqAJWI2ajnR4PCS5/UqCquDw2hoO2TpqSx7wVQ
9K2PQSe1nD+p9S10tY4wzMfqW+jxiZjm0ukGGfSlW65UEWWk4S0Zb0HZtrdeimmr
UkRAxdmYmXGO4NkdipR+MJhswUbkMld06/cxDqKaWWZTRg/MfJ1LheTNnVgA8uLY
Rc6otiPNAIfm/zD2alOM6TxrvrQaz8zavZEE7mDijBnneNPZ4bW8xMdeP09VL3Ce
fy7bKO+DegfRT3ZQyzbpANs6EzhFziWACI/PHVWnX5a7euArt4Eak4HfhEjMjeVO
IAyMeARKs8ObtzYnqEcMD2YkhyVb9guu4dAKlxvgJqHZY5cSHx2tGtRUiXNyuHA7
cnT/6xBzPqrGf5Vq5YX6MpVuNIaT+VJiphxkSir6PUP9Ax/Q3KoZFiWJ+B9jbGK0
dPQkyf1hOoH24RkYPrDrum/B/vULva+5E/D8+9VBnUzvi4reDG0W68++FTBYCT/2
PZ+mqOLNi/LI4s9wOCSVq5jpgIOmLQZxOGA4MNzkhX+yI9dneyGBAl9uDKa7EWRe
WbWDhKCMBSMiBZ62TLiPuQyqfk4AR+F3XO4xFcF+UnYGWK4cuMLhlXvOfxiqa7PO
sWa61Xk9M+VsyT3dpNo1l87/CgjXQsoWceQW3+vrZxhRXaAfnB+l8rIjNVj76bqX
iIP1kyA9UUBoU8yhRS+DtLWSMkXCsSYQdMsHt0GeBGCLqLQQz3cHKtOi+iPzPQ0z
m9cmgWiOI6m+J8opbtz6SMywBb4YUlxjtxJqP1FUirap3Cg+enejDEuHB2fPomIc
ZOzkyCL6sHuyInf2qoAmQQp3wEl8dWg7/72Uv79GcuC+z9F3WXbWjANW44d0QDTN
wAL2jxDBL6J2P2qaCbBn1KwzE5nkx3ZlU5gYXUspC05YivD3u9crlGckkSHmZZM/
ENtNdzmWCwxAk3iOm6DveIHNOa1ZdHvir1FaYMLu3Y022Jg2Nsja4FBSjbCTk1AT
E3Uyb8rkMWGL1cT6dzNPwdaswPtazEPGMSDcVyBJT9ZomfQ67mX6IOWNb4pYIgq6
/kVJGbtejVl0F/KXTlUwAUwy8Yrh9r0tE/muUVS3wISssqsNpU9uOne02C9Wx02z
CIV03StmzLf6F6xHcgWmCHiB1FdFUKNEJKDHrj0CxMRhX1/smMIlPdNflHRs4nmt
03GHkXPsXIjbguyzIL7rUJtsB1BAP+BmkYqaCXDpzlyXXJE2ZPX/1ub4FF3/1lwd
uToHlte0I8vyQgupjJh69Up7PvALLBe3KvR5nQqpXFeiRujUY69uBb9EBHtsyPzd
ASZx1BM9MpWtMzIdeiHV4zmgACbHxKJ74UXtpRD9+r/lw54JO2CDPKNgud/RAkbr
2ZCjWegWXe1gUwOF1vTKeh3lvCMemlLFMx74v4jQVxZwDsMzjUTxwaORSet46cX+
VRjS2g3yg32q62CKmeLkoVcAC0zohKLalc5c0ldGqqsU/4NkxIprMGLGn1r4IvGz
QyL7H24JY3iLAyz0He9fgNI8O4p2fQioDTz69FWW8bhrmiVavOxe73XdnXo249ow
3Wt8TQ6phg4IuoZ3EKQSOrlPc8b1ibc8lmAtrS/cf8KA205Ytod4FhGwVQZa0Mlh
3rp3JpnFDO01H/nADnn/KYqL1yiTOZyPHrLKXbd/4VheNFeZ1jFgosZywI/AXUXM
1ui4yXek96RUY4ObFlje+dXIHAb9RJ7CJh2fvqOebPoU+zPAn5LMeS1xiCdRX5mq
rKbcufhKW5JCWgNiWoN696kHuvZ3RxSt4LhAKkxu04zgWD0zJmIUEMaSlMGZjy2T
KHAe+yDtk4tE4MTcMRMz8+xgp/KmqiGQhsKyNwuRhcDz1qy4ISkCkC8JWJeIgTQa
zxYk21H1KHF5R9tzHsDJyzVXjwePCW1/9zKT2jMGlGXQmG4ksLWvzPmOxD6DhfqE
CH1Fvy8NPZwXrHEpRrg+LestMNInRxsuRgFZ/vTakwoJ6rTzYBU9VP1ao4bXSJGl
Iwbkvwh3fzj7U7CrqUOIl1TVXB2CBNvUE5qWw8/Gegf81A2Q42dZUDDUYzq3RLO5
wB7heR9NEcF/THGAhOPPmkKrN3kDWYMSA2ERb3dxFZgMqu4Oh53vjwNIJMzvXSow
MSlqr6b8gCvF7bjVUw3Tr2elMVUxsZfeUDxcSYk/RgUEsPyXgO7FC8EyEHUzLt0z
sKwbkR5KT1WBA8Y7WKoBOMSVPSJbbjRoKAy7ueMq+oXIqy0/Q33Um0iP2I2agCjq
mO1H4numNTXrKtLcZFNUprOBAks2oo0C1Gs98HDc38EEbKqwt/OaZu+1wIqLYBci
m4DXhAho743bm2fywd88EphUvCoCEdQROZWbCkU3RwPW5R2MBJuuycOs+D35jBog
49/DUAP7Ia45xwWXuahRzQYh7fFOAcHH1lveRL0Qz6pYQBJbRZR2kPvKPlaua/aK
ZPNeT0R6LOUbg2yYPF/D78pPN5qfD1c0/XMYMJwSskYW0aE4AR16K9ux9Q3yom/O
VmV4CrAm3trmFYlG/a0iq1K26kZFEuYvKgYP88AA7fbh8NF4iu8ePQJQ3NYuPKgS
NNDcTD7oMo6PDiscbNtvgTqDgjV3U50nLeumVLIro+eSOAfsJDH2hsXpRzI0LyQP
9WHPbkLnoGpLfupuNF5G3e2V/osSsbvF8kxt6K/xsT2glSRpN4VkqfCQiuk06/pJ
T/JI6uiJSBoTM1HDb421e8jk0nUNsqn/xSGiprNKUOxuVSzbx2rZJH9hRfm7qfja
TREbCIyiF0ACqXvCxD8ivPaHrnJgV95QbT29Tqe4UzAfDyzFmksNgj6Yta8/n2OV
/npPt/FRgsAaZ1ePveUMwfRMQowGQZhCUQvMGjDMcXHVTfsZTu98k3LJOSDVSQ5E
z7iUpUaPdvQlfqspZ9+cI8FkBKGBd37UO8Sc3GOYOe8lEtszak6AD1pMF9NVO693
jhNFoBZZepP3KP4x9JpfwS16R6rQZeV6oBnnk2V7OavQyQuh37vMbTc6ej90dn2N
lQETgCCdgOef/Fp0d3sF14Yj6j3en+h34k1DIQgtZtZ9gxxogKOoGsIzHmZV9DM+
4ex3Ji++1xElnioEJ16Wdy7DkPntNlqQxJeezYcRG4EPq9X58ioMoYnhNn1vzIma
G3Ozv5Frj6+YPKYYX1N/MXTyITJVowF5TxdyCxx0j+yMGIZNfjCOwthHsfcd5Nbk
PNSsGDURcB7jmG6fNiNHF+xSUWLH/r8fsuIcRnIaLEYxF/10f49Yd+dl/Pry0jgd
VmbB9Ra6AZR1s7BLktS3e+zHAqJqnexk2lKIMhgFN3eoKfXv+Hc0FNCyR0Cjx3hK
rhHtjPNVrvMIovjxf1pooB5rwg8yFPAeckWi8rkI7cXTvC94EeMyPayRGNutzAH4
WEnaQBz/D1+TRIzl1dyB2YT6S57Y7ib6Os5Wo+X+tiWjJtd/Dq5AHZDiwdzAIfJx
nwNg8jms99pxxuSLJuwtZlRcL/5jdQMbEmRsjaf+z8Xseph7+F5EUH/apwP9vipZ
cok8nFDyglwb4dEdRPgt/1e09U0G9lWoOyLGIj1840ShRmFVSUUdLES5IoKcHbnh
xadpQAmyLh41g/tCNqknZVRnW8WaLprpT1r+3S/lAF0zLRBPTI544yXX1RyY1/28
I1fO/IiEF15tFWx8k2pZ5UmRiPHsEbEuUgUECRqddaStTcsKDY/Shuu04rRj0Yld
oPwhKq/HzYmxp9OcI3mJcyuO2mLIO3r/NXydZDsV09TfkhQjiVQ5QdO8CpnkRt9O
dFq/WqyGWN2EdvjTkwpYTK26oQ4adiHJAKWZmICF2OyM7zz8FLcpnfsIJRvu3nqo
4U16+N/tRK2YrPNm5bhZAG6G3gKQP01KfXSxkIPcenca8wZrRHie5vWps5HAbVfS
kCvhk+EwkRMlFCf8QsVF37G1HG7/gLjqudHfMR+0a0h4JPGYlqF8r8dPMYRqNFmV
7g5PoCa2Md3ckSQNRIZS7RMGy7/MHF8AWBdRJZfYrqxiagdHe2KIREBmdzIqK8Mw
PNeKuIdhvkAVNPtEx9wfzExJ821b2S6UafIze6epOJt1yeqJSdKMwNq3upq+Kak8
LU27y3671R5hmLUvzSybgIIV85NNQJSHozNQFxiMHpmR72FfrQTFeI1MmcZZn8F+
qpJCO7MnU3JWI3xNT0E5fgFAZcpCddxRWmGMx9s9Tc/BKo7tyLwHJYkcGJGhChWi
y5ExMlmAhFnKlmqMALkoRtmeXt3u3cKEIveTp67bNl2MXPdsVV7cGO0L9fyeS5Yf
FbNp3HZaP/Z9SWHg1B052rzcT/BeCg+FPRdOYd0VmiBSoVoJfnqf8YP6RJZHrS9D
VRDmAS/5/KhM7B4cLiP3ZUujUobhBxLTmxuDzSUFvItkqdPBYA+CzO5ouDTCLIDA
6Bj/i+8DNmNACjho1D2P/IHhRaXIZm68ce8sxwpthaFoSvXNrA4fdeAtEoB1w7sH
5tCsSSl/oeeqSHX5wJdoTQlBXPO9YT5m+JzrDuFC6EQQf3rVycWvPxMFDo+cmBaW
csqyPH0186YqY//hs5ZagDoDBlh2x6S/3XM+sDF98ysaB4DLEPHUxQJBkJ9VCvdS
4lYzU1ETCxma7CyLj81Z9fJa17oLDlCc5kMhuWYZeBXINozIOt9btUj9+xhJ80I6
L6VArtdCmADPsdiIrXsME51/RZVrNdFzlZJXI1ikjLm1U6dXspBdQcHoKFBFVWFd
ME2NirwbS2Yo+KeKe6g83qJN1dHbNmaZqMWe9FILiv15dq+AiMSqB5aC/9JVkhFG
rIyoWzlM6aNemGdjJKK2URX6Tt3KDannvwefJiDO9swF34w1ufpDyspa8klhJ2jk
C8/znmPKsBTels1GcQ+4haSL02HEZkkAqPlJfaC4XCtJyjFbzgNlx8x/tbZU9elZ
9Jlnebac0B8sDWZjBYpzi60+yweLysZbIJxn6re9zBchYXQi20XSlYfHUJl16rhB
eiY2OPaf6c5UQk2TAJQw9oPfRsSk4aKHUpDvk37+lwpp/07JsjgbszaKt8soXw4r
Bh2po3IzHK9vkFOg0SLU1M/kju2tpBw5cYdC01ljX4sh+CuATf6D261Ns3J3zgR8
uLBDgGoc8ueAgkKxB/6W1GowW+KAkK6Wsy/T2IqR5jHAd2UraKmUHz/CvU3TPb7I
1KObm7Y2KCahAjAH+ckzOxyLS4RoZAWrdBeQgBlZwqWgqIqrHJCBiqQm9Fj2IxDq
N34jXl8srKxTHKKsg0C00OIRUb8pRsoDAeJxC4KKBjaFt18lBfEaN7VSDx66m06T
Gf0RyM15hvmvwjVJOzmTu5A2pR0ferHOxFWRUiKcDtQzrr5x6GL8ednkfJV3Ub05
rR9GSCqtQLCX2ENEV8enlPOt6A51lQ31nc/Mp/GegW8OrEBqjjkw9WuFiPk79/rq
OGyBsrK+6B2TetpaTpR7BsHP2gXi3PBu058UF34d44oKDS5DiS79wiXhYrXaQjdH
sgY1THQa5wPi/CiBW23xZQP2L/tI1si5Uq0koVGuznWZ+Lw6ska7umgvDmSPevKX
P6reRu0tFZp1gCIGt19pkLAwckAbqzrnpj9mhB2Jk9npbFkBIlkIzJgHiPVj2tAh
rx3Mu49cHzLZe2PvNIQZZceTlLYkXcrQDg9TP7tZn+zo9mbUnTuhnu+SpS3Fq43x
qOfq4ajRg1JP0GIh48+1bVyLT/eVuy1g9GSR3Z80YWk1PpeJmp4GJeeOK/6wi0kf
ejCRQ/L7EIfj6D6DJdJfLP1rAm5gHjH1TVLI+1Nso2mtGvoAzpS2xBq8d7lg+p+k
9/mS6Qyi9Ibo/Wf/tT0fal39+T1NkDQ3CgLKldKzvT7ry7NJe+oaGqkNveiHzAEc
foiRUX8e6GZN6uKxU+ftgY1wGKaB1AEJ2qn42mLX6WvTtrESmMLrg3LQOzX36amV
lIeF+6Oqg80VqsPDrkuDtbi9XB5bxEZotAqZPsZ+ik7p+S/MWoQEIFiDo/+1CiqN
PciSznwlWBf5yVVWJ3xsB93gS/LkUGdqG5Cye2THSy5A1hrh8mnYT4EG4vXGTL8k
UR5fS8mDkNozr4cuDLJYSQp9Nx8gsHpKV73dxa/1nmVNLnnesJ2kPKRs7Uxrosrd
lIb7wtIr7DieIJpcjv90Kll6GswGUPD4wk8Ab4VVsAzVIKVo6/KjzoeN+Q6RLT6m
9YOsWYW5dIo7wJX64NrDrOywklsy8UEvJ44if4PIpT/AOUfqZgBe3IXpOYUu9JcJ
PzbAJ0vpR91D23Y8wGzzDkoZx8cNMFgt+FQIymiOOuKMPcbF/uj4d8l4QAirK937
Cn163ksk3oBPOAs8d7832VmJy3z4PnXfNnxcVqwzbe6upwSTrnsfh8A1h5z+zFQg
fGGkxsTevkqdZA6buU5pkoYB+rTBnBlO1JXplZzIvKMFeCwvaWFkDGVrE2Nc/HCn
8VFzJ44zjDR/xEYLH8wKW3+zGxnyQbYi3TyraGPrNbzbxHtf0FUZlFaD2zRcTB/G
ahYlT4HQT7rGu+mCcgZex9iccr6jxKM6nk14V0gDhjEM5SKHIAk7+uGs0VS0Di3O
unJeyiPdP7yu843YlI6dx7dMkzq3uKClu57CgoyPyrBgk73qoDqorSZKf1CBojV3
ng36GQnQQfBIZbScKwkcz0ggIrWI1XrhTDjwSXUuOznsubljUcv0TnuFyIrJ77FJ
KN00LJmsO5t83bhMxztXAvBsFpH8rteZz9ioaElkOu0I2L2Kiny6lVxBFmd7vNRh
yCBhNhACV2Hvo2XIRghTQncp+A+y5uzLv3/95N1hrdvSl+mOIoqZjMIhnZetRWd9
ldI9phd2+yaiJwfpqsoz5MlPwqiF3z8HpKF3e+3eS2/OpNK2esK9dAVLITk1yEbl
bEEKXL8MDB0NtcCnwa/+uJVA9iyTEHNBiDSmJvMTfjVWQFWP2Z2B6CzSNZDSdHxP
hjbZRL82jEGKuoheIbFhFRn5YpnR2eDEM8BzKMJ5ZDLCe1Z+RXLP6qqNapwCN2n5
Ze3YpUTDGqRnKbZ4WhVH4fNWotkp/jzLtHHoxDz3pPcdu+OZuTn/AcGoFnJJVdzR
Iww9ddjSYlYHn7Auu6AckNZK622mZv9It2w1keNyZvBGaEpYVRimlmORoZxRG/TX
Si8eXXciaf2ttGjuHJ6fGJZy5GValosQtLKOWpPTTekfRRhg/R8yoAJFwJvYXahQ
oI7YqZGmC9YP6qPwIEpZJLdxTwK6VaWeR6LkI9w5S/y1Yufdozxf8KWlad79rGI4
ThjrMynF3KZDscrRde3wpWsTK+T519O0eFfdHnPvhzWQhw9M83W55BblanKBgX8l
vFMlwHhG6WE43rYAPTwc35aog+bsl69KL9Ixni9eO8AMhx6SBDn3sDXRy3TYG3JI
V/p9zwqLYkPmqw6n6gqGAdmunLZfk7WJ8GzadL1WCfwkOCzEdoT1X+Mfl8zTkPit
jhQDGPfyGwzZzLubc+xRfzXrFdicmaeuMi35ensdwMmNqQ4AHZoq1ehCpfyaIS7H
1YRoAlyevOuBx70kZ3HDwLWWlr0GIrXhUV8ftxQmEbzHSeWOqCIw09f1gJV0+dG0
j5/t3dRFk6GJ8tOwWsKUrsEP6dZtYCup3HajAn3LX/iyhhcD0Djkr3Ofi3aFdMcX
VRDHDD/3rg3fKO3OXt2TR5TbBAZY+tFDAoolvZoRsICVzstZyKkPnghkyZWlAM54
zfnKGP1ntX9p14mbJmMeoFgRBPl0/PC5bFwJi0hKOE7wkdPGZsRAYHNrplFvLonK
I8SbS/yoRluJJa3zHTFOqVgP1YEHxq1sx5aaBEcK1jvilLyZoX9sD7ZcQTla8S0I
bEDFLkOFTFUDR2Pfvo8JhDw1QmIblc0NbgYgBeH1TaErLirafH4Q2JyVSK0WX3EY
gg3g9iuMm8BOABu30pr+ytwoT7ZjpwpK2cIV6MisoBruOoPEA9UIOGrVUthPGTOJ
BFmKuAeC94QrrXTFiuUqZYOt/fkrX0tRCxcdUnQKx2Do9q+3jrE2RQALI9o04NAv
X9Mx/ABAsPb0ugGLUzlFN/WXX4FLoMxym66VC+y5l/O8nduyiPXykEu6mJ8iEGRY
/Yhwkd9AB5I4lrwkAGa1h8NBZ41pSdv3lysBOmiZn+MBqPGfb7F0UipnWedoS/fE
K36sDQiFFdqfpUsMuizZQHXHJJD8b/snEsYU9k5yWKxYBkuvvxARysEpT1hrcPQ9
J8eRBU9rGDk0qPMHOvRDj8u6DOa0EUP9W5a2GAdBFE1SM3tQdLOxpsczDaS6ajNl
ANzckiNqTFpo2baOyF/8GUfOQV+Q4Izbf3ZIKf2fH9Utnweo+jhELlURbgM+XF2z
ORKM0L8/1P3KUBjNBnTwmAxhUZRCn7yPx7uZDlhR3vcSks2h/oTExnL/U7PmY/sg
3rDO+Deqgn3/HvZT9cHHLGU1eXd98oWR+tTdSVb6bOlwinS56fISow5f+sK27pr/
I06hULKmfjAuV65AAc52xq8W2iA9yHGsKXnG3Ak8S0Yp6obvXCUFwnQeNM4m8/q/
RG9wZJLtGPtUVOffXGdFnpsBumj+HE07CyeSkDlNHrtyQtBSA7p4bJzo0v9FIthM
Ijz/hqHPKKpAVBgEgtoKDATHksR16Zjtb/MHaoRmq/dmyeFB1kTS+eUdMNxX8FiI
pi8wCV25raF+XxGqqrvsPKMOPfctEXQicFKM6vw1Qd/iLydNS7a5iv653wUX2jxy
/rkaFLU317Ul4d0tg7LsLggtzUsdy5zW/7w/BBdxCwFsniu+Y2leTJfGr2XYPG7y
3fLQu8bSf9RBEItidOQagy3Isr2JSkejr3Ilp36Mob7h/AiOG17tkWbCFodlP8wH
5vRwQORaYz4/YtimG0JuIV6vzijXMdKlMlHR7O5eP4damF/sR/dZlyO2IdWYeQ9e
o0q+demH7oQHL/J7I1X454oirxhOw5HBywJ2WrcFQe3/b4+q43j5sNPUPlz4f1Jy
HYYgdovhoeQzMYSajt8X+DbZyDM9RyYesLWRnqBFMd4fUYJGvTyN86EVr9SrOM4i
Lu4BUn4DVSGK3Ky/Itp7x22IZBFW6WG73HQvuCWx45SXoG63sYOKNXAPRZ++5V4O
oYDrQptaD4zXos0932qMdJMyW5RfKExvfYPmmm2r9b/nzYR0ict/c0uiUIJsJxL8
JNQSzgaDllkDFV81+IzaY/OTyr6hqvVt9E6ibtLQzq9Fh91Qt91ySM7IeSlL/YdH
wM+xOxSBTl28FIgCrdyOVB48IY9JSdH7w0ovd5smd8SetFtOCd5qkibsvaxTKCxA
kLwZFUo/t3JfB+6Bnxd2MoGK6xqP2ZUvXpMAZji8uq4FQomzbuaHFiu5auDhtx5A
oihnDcDN6m3xFZqrb4I0+f5CnHnCniAkOBXSLQuI7VWKl69N2U1RydWdsbbze7E+
upqh+2JtuLKX6XlBt+zRs/urQdeGejMm+wBQsh/qtqap3rwpZmH0ZBfpdV7Y/YdF
DVkJKSGoux2ruPCiX5WGQ2EdGhQRJkrql4MeiGTL+eUQSs1a+IV9yZAinUjib5BT
EEuTiHy4BkKuXwn3Aji9Hunv8FgjC6VMzE9bB6XrQqrg9zTSZDxE0Ut8Jdv0QkqT
K3U2h8TqY87hdVfTvVmqEJO5oCanfxi0YsfPkHdXNTvgbYJ2UpqXyXNhYW3pvrjj
9YywsmAg30mhv/+9Ix4Ru7e4qYkW8ebTJWItQjmvTLHnMPswDSCkhAeFW1pR6N2D
Nu5bJLgl4E+JQ5++HKHkb+xZu8hskviqI00+3iCghjMX3Wpb4JAt4EcE2WmNHy2I
Mj/7DpVsJ3zmb2kalJ8dkgpaaGpoaqDm2T8UgufgFICT0eyOeHNoVZ4TE7emDRF0
VHJXpdyek5qpT5NizMuE8++Aafj7Z2XVaSD80HcJFMrdaTh1lS4DbymkrMkOQ93u
Q0GPVEUy8Oh0LF7X67Vry0gzWWpDdewJiV2bBZmfYGgukJL9+j5Ufn0dbkjoAmmy
mZRzYeNSJgVASJPLd4s332mxBq+CF2O8s6KWp9NHQkmFNU+qp/I9nJebYoOw5aqh
gJTUylv+scRC0zm3vx77OVpFUdCFtn0m4UQGy5RC0vX9vA/0x/Q5dXhhLy8LMMZY
PrlHa3dzrJFcMgocdCj/Vo+MiGmzVrc4Itvt97uxTww1a4/7Equ83RwUZKZtPe+T
5Y3XkQxz8fw6IuU6WqyC8FY4tkidTtHGR1v2sQI4AoGe/InMEnl0R4VbQFbX231M
+U60htOSeHm2qkZiLL8O00TUPOWmRRhTzbsxA0dDXfUXxhS/XcMdft0YZuzibbFO
gC5NtpBbarXPm56nDqMdEh4gDnuvT3WdPbRdm/xNXsTaFNQwS++9s46TSeHklSCe
hBg2oJ/IVP89ajBuyVjvGwKakjXSiH3UiFhriCuXtwrUIqFvoKDMdMCMgcG9r/+O
7g4kKljcxezTh/GgEa5y3eGBecHQ4bXIFHMQCwzetLHik6mDE6zNvLFfKvkwNjgS
jNc+p3OQDM4v3toHYosDkmitnDrmaa2EeSG4iImo54b49NNFsbAo8Gnc44Nojjmp
VCn/7HXwXb+k0LBigG2gSk6lIW1UQtPJWwli0IsSm2tYRIqwcyKpwvc7oak0Uk6T
kU7cw0YjvmSM3rM2PmJZJRvbd87DeR+I88siaqVjBgDeIPY+5t9yVGdhgdnNAyUn
leXVT7zBEYx8ny1dCM1NALWRTBwpRu+uBmmaXDCFRShPrTmPzKSlT5TPK5Tc/xGF
CGcVBpnRsxZphQYpx2iYoyg+ajok7isXUc7S8ceBOnpwQwPDqNMAhaNtxDe7bGkN
A2rFn9Lq9oH/Yw4VE00+DjRKnqHeLPYXGxpIHcGdDNgOimaBqeGWHjmLbuHaWf53
67f0ZhL1+H300YoOAZ9lFV0HnzuF4jLx0dH5DudmFoqF/b8+7/CDfOULu/ETu9p3
vTNOPj6pgEJY7PZNtjsCWLuYUqx2zV59iE7xvfg9754vJM6cqJPWSdGvgaNa2Ocy
ze3erz9bHzTvaKABMK5LayGv2/1Wzth1Bf/kHCeVxi/r//7W/LVYQH4q3wUF5oJc
PPRQWayo/A415LiOkxlNPOBfUL6smnq0PEj5ZxizZhfilsi4LSnvhMefJIqtjpJK
4NQUZdL9qywzAO2Ew9bGwwZLvjgpjQmO7zU59/lfVFEhsQWm9VPMvBcQhtwoapZL
EuxiJrjwueziZKCJIizx+3Z5xyLkBXikPHOX6W/KYI4ThMq9/jAVB8OfCsDAWaUQ
CI+1n0BMMPybFTcEJUHJTa2GfgmbFk203pElG/8ye196IrwatR+lqiw3Psl7P6po
fXoxC3HOAwCU05ABaomL9x00HhzOhNPt/UwoposRN9/SWVbY9VZZ9ol6FBXrpkPh
ZmO5W56XHl1O2Z8KuMW1TfYEobzWHCtgDhjOs4rOEfc1HaL5kW8QhAvgUbMt9DLN
7/RjcDaNyPV96dSHH6jAmzaUTkwXVzBpMDJ4TDeKU75InI+z9NhUXKcDqzXH1dos
5OzWoxlcueZ9jFMXkgZx0QLvWP0TKiyTuIq0qbsTyEL9SqaR8T5KmeNroemsdKQq
dFqHV9pu1mDmVCKxCM6QeGUU72eF3ifxEYY5AjhX48cbthfrgfIBcgtcGqeqN/pq
IxYO+qifFp2CiJcyBa3KaRlsok/5iMUatfYPuhbYQW8J3HS5po8/IEiBhLuiN3EL
iLcBqYK9a7DmQFz9/P8fcmvyRS7WZjCxHgwERD1/fHgbaGh5nyX0kxTM73EYaaiW
awwHyZc+duOlDpZsRt55WRKv9VFGL3rdMdtyHoZRUi/kJzvqiF9nqXurOCZHPb0Z
ESDqYOcYkqX7oSTOrC7Pt7NbyOyWjcjBpTaaM2nDv/gXlip/fs1W5vyURxdx4OlI
hleOCbXTUZeZd/9L+BwUGPZPyJkucLkZ1rbtHn2bF7sJ7DGeR7ZgnAP3r1TnfEpn
csq2Kk1dOB4H/yLg7U7Xj0wRkztlfco7yqr3aOen2v/GHIsb3byJDf9dkLZ1q4I1
fcez7Nm59wquglEkX2qp8fq5/SfGzehzYJmyfW45eQYIWHNHmYpEzoKfEHZ0Mv+x
JLLcKn4oGFDsjyLCJXmPAhc+isprPmKlXO+noMQOqhz+QjzGwWaQ34M250wwupCD
I+ZLO06gyVO6ap+hTx6RvdpFz5IezLwl4OWGDSGctS877lFcrcCHbzKvZek5UoUQ
jfEJGQ1zqY9vVlqbGYqAlVQOKQnEiDcVwCgduPMN1q+pq4szV9W283lKuKnrjMDk
uK/KwhZtPUGhdrMqE+GTY+ZbooKGxxZipWsasZ1a1yhrgtcxOcx9gi+ZAp3ooySf
tjNDGEQAJ/bqjpqDusepxOJX+3tD64GbjBKDk85qqHEpzFULuhV+zS9GzWDYo6Jc
dstVixP/q6INlKmERK1beK6jl9JnKH81s7DX9DSxHIbpN6+RS/eOHKtQT+x2gnYg
Og6uONRAlLMwyNpLio2dOneZbVyhaeA0b2IKW2t0WqnijorolONUEFcc+oxb5eve
jJdbEw/lwaWOgUoGp1dHA9EIh7VjVU97A5JEQbd8M8KmQqZU3DhIQsfbqW8AiYCt
vly7+spX9GXM5+yH2dk5Uw851sLZINShLSvL4CjMsv187bIKQVSzGUZBeeFgTxax
YcbptXSlePY3T0uDPngYOTmXc4HuOe70v8gaxT4LVUpmKndK4Wz5aqYOL6F2y82Q
1y/awyO6UNqBaNHkaZuVGbAURyOzNaT97TkLKe7FTCkjkQ3nhpolprihkJSuETlt
B79dwXCD219w3PnyH239DrjwF9oOzWopVcOxwY9ttGAq+enfvdn3LxaMrtx4iXtx
fcf2S4NDsdoX3n4/Gh23cyY+d+qS3jhhz/A0mHKttQohQXuz+8kU/KsqV6ayvvmw
wn8GovJ6r084V9i+7qlXlKRs5ueZZ9rv5IW6IjVOC0ERozgYJSouvQJ42Xa6Yp/b
LahgSAONe+Eaonoo6JlgyWIda+QGp5htjaHRMSjaoJBl7rXIdkV6+ARkY5f9zTek
1jTr9NaxmGLP9dIYodfmvOT3RtwVn0jzsqrNmgFgqp163DW4uAw91rn92imf08sE
JI060LPiEJc26KaMdaso0DsqMc+E0XUsUBjGOtcHd93Y75b9D2YWU+vsFwD/gBZA
y0I1BoD4FJiTeTPegzd/nk4wtFHCduRAdXwRPCsv6UXfzPj5dKgEuBdJuM5gtzQT
a5aec9LURaajnzIKnC9a2SA7FP2OylEHdDToCaoMnQ62tlwMOcQjSmHlHTBf4Fkf
kHyK7gol9JHZGmO7yv1qnNRZRZmFw5xe1sjwtpZlCyE49+3E2ZIpugaFpQO6XJ4G
AorIiHQgyGwORD72ASJt69fjk7Spq5G1auiKmFH89xbh04VLDGIuefOiE/NC80tr
W9w4Z4QxHmx7+8xUdal+jCWfFPXBskWRfcdxvxK52IGrWQBpDHDYYFh46kDLKM04
3tvBudlIKHOXAA0FsBIjxvN+iCM8Mq2XDmLKU71xKBq8AR7oWTgavMsrCzyQqzQ2
XZ38QMqIOhzmH/QpAwkm6fP4NUukp6ausrdo0+nR3ThDsv+3vvd+gIauTfH2rbNq
/SFPEfdCC4NMkG1vLV9owHuQAGY+h70sxTlW2Xh+utLseLD2V/Ud14tl4jmqW3RB
RuV7NpFROF84YRfbcBg3mSoHbC2g72/Gx3046LJaEO7R7HuvK1uLRfBFkBg42UO4
X7XyJc0ZDr0MAkVP+ZygQWQNxQcVu6zXQ/eW0eCDGfNKdgCOyHuHw/6Jm8+wgBcW
eUh203pVTpdZMlzbikBlpC9PqjH9q3nHyDDyB00OMx4FhveasR/E6XDKVa47E19a
c2ZIFClGTJirGY/Y9hZjE446N0KAxuWf4l9r6JMGdzJM9EMzG6HQQSztxVkYGMMf
Rdo7ouP6n7tL9VVH8Z/KSYnpwYeYzvfp8hjQ7RNo5LhkgMKArbQ2OCgvBcC2FUoI
1tqgtorSbsw4SqZc0VcYmpY90teZwyk111CwG9ZFmshDrAEdLbby6JAgGX6gaBgZ
rmHdmjs7wffi8ushGGdr5alIVnah+e1+ACbtsgREzw73e0N4oVeniA7FV05oH9hs
oxVQmZ4QFhZTenf79SieoA0DHoYCLEaoqzWG/gbKQYWnC1puks7Unb2zR9itrWJX
j6ra/pGGq+aHN6l9IarzcsWON2mCpQ3w9ocFnN+aI/JThvZ9m7PVJa+lq9iLUnSt
/2ok+z3bnHxj4b8EXW4P9wrQKgJtsqCZ9Ikdz0uOmxzRf9Sx1KH5f1iLjaRV3jTG
tUeWzS2CiGhMvsS4iYv5LtXvD0kQEfRRuGFVWV/it5PgALVvhhsUAL2SnUGRedHr
17/dAchaWt1WM2ie0BnaOhHVLnM10RdcemLt0Y6JPwaXG3iGdsKRFlMY6a+jdynK
AzLOlnFc5wV7xSb4UjIzBwtUN7VNF7vTdccIO0p2GyPwi54zfNKa+TLPYG9yYTH+
15ljzFks2aXImjUD1qVhq6o5yCr59VIEM4Vx5va+uF8In7lwNkCH2ouEARyOHHxM
GGMqENNTYLDKhYzPZIUnIw7m0B3wzh+9tf3OBOYJtapBxLqbPBRjL0c4QHX+Qyr1
ouGLBFalEVZYWrPRa/Ks822zhSqdFw7n8UA4v1xLP+zhWh8FD7DnjcQ0Gl+exv6g
ejbrr3k2SmxBc2QHb90fTJT1RLsaza8uSDOz8PB0TH4EeONJH7aghNbrnM0OAKWn
u5Un3tAbDP6llgo7nOn//ifXwBDRzrAUpjlbJPlDVkEGrRsUueb3n8dzphV//gnJ
FnF1/3a01WhD7LtRLivg55PLiWbNrcuPNzsOZxZ/dXKBcm94ujJhVF+ZnYFi6k6I
2dpunGLew9R0qmlvMa6vc5oP7MIQx7XGI5xj3l4NZ7vs4O4wJ/rTamEWhekLbpst
0qDLHGsbjftpeUk2PAyfTSWYrIr6NzcZgnd4oLNCXa21jhdXLNkp2KYKCFdMvW8k
Kk36uyrS8rdh1DE1vX+13reXX7qtKRkLxow/MaucP3HR9O4XcourcpbQ7dbiBO5e
GuwYdkl20j1srYTDF8Xpu5+xKkupkCItJkkFR2CZ0ih79IKjvcSc0nbtlkl3YdBC
DwksP/+A5kf/x8pfSZ4sIMfC02gIUI9gTWt1868dt9c3GaMwc8d6j15sArDK04Sv
CqcjHG69/rKXNYW3xF7eJ5MIORQJv1KGB3qPZsjs0PzH9RvLWlJ3J/98twgw8SEo
nQnLbPT1ffBd3i/HVJG+yMuQaelEK3kTtt6A9PhMFhdpJhpezI3kvx7ardGFtpt9
bpIHei4RHccfl2ZmmWDAIXYkny9qFjbvDlA/Xq4o4AIHzOiDqp4wlB8SKJduOOaX
3JDkujbGDevVuqseIf8Ad5RFlkiBgLAK4k3OkOkhkU9+9IZI5/eykFrCevPzIfPT
B5Hsgpt31nZXIt5Oz4CzsNCy747KfoAI8/3jMgBgOZpS4i9lObHAZqiS8xBSpJa/
43Y4eprSfL1QVGilox+CEn/tibD6NSH4esLXKw1A7nJKaTWzavSS1p/EdRTQwzMo
tG5sH2MttTvin2MeH0qFjmyzZON8vUmFWTz40ZtcKlJB9Ir4Z6kqXZpM63D7dhfs
6vDjYoCZttT/QQKHbgW1KI6UMNcWrWs2IKMzrC3I7fuRQ42bW7vJKCx5Ee1IIL5P
Jz21KX/jTKu/zr/pI02P+h7cn76MgDkmEVnZtDN3/RIP1dYwNdJRwMER9SQZxFHk
jyRymBX+1RN5BCXdM/AxU1cKski3K+yixuOy0Ey4llMtn1lXS5PXQrbhfRh5ub7d
YmpVcTha9zJ/psXAFhhNSVRvnap0c4ZFz95xG3T9AWOesR1HGnRGeotBUHaVAQJU
Ny/cjlg6jJqwTCdVmc0H3Mg1uqu0KJ3rj4koNLNX9NDDWcWgpQdOTtO87EzkKAfx
UvntFem/YPgV5w52JhNMIwHDN07U7MOaVdBmHGCeCh/jYkMKHX20WS0gmV0mSL85
0QWVVkTokp8W80osqnHPsjTkP8RzwKsmune9mD50kS6ruczcHk2HSBMQs8dR34W0
wypO4oOkkn6T5xjsG1Af5EqobHIIVZADYaaF2lukME6fk+Iwod9QMZd3gdJDOGNS
nWODkfIN8JT2urr0jg/z7izX0EW944+GMKeYj99nkXsV9AIhJeJOeVbWjcRL4VJi
HmPWum5+p/TA/rPKEznUWxSN46N0FvdNAsHBSEAQPF0K9WjHasfNWEcvYu7BXZeJ
ubhdXC+dcKkuqyFYBcV3Ik3DyYe/f/oyxKWlvy9dxbABqtzG2EboP7kBMoLbvKrW
MAP61iOIuk7mR55bXLHk0Y4YJIvAaneHNly8J6jUS8Tde2t1feWJ08rPa7/ZHxiA
hMTTTyc6NMiTdKm/6bqIdgoJ3ywZbuvTe24NtbMAnQ2h9UAUEghva44cPbR1PbTb
v7OUclEyOldxNvtZpllamnG2r+JoNkyNpAzgfpDNBRAvG7pg3KHWeXnpj7kM4QEp
n+WCHQDzYNUHe6KnrNE34C7C6D48ft8WFy/vKR85l5+KJ6A6XvcKXL0n3N0dcfBT
CnjlNk5NL1bkUR5D3LVda8Tfsu3B4e5HslJE8fSiog975S8W4SywYb2/R4cXWkj2
b39iNbruhuLRnW+GJx7bcUOK5CqhGSk9Ot66seAhUEgHeZleRUDCklfwcH98ui30
EMBObrJVPcgYDnKzEhA/IYTKAr6ImDeJZ0SrBgF6gkQdo+SNOMxyhbeqK9zC9Iue
Sppzn/4gnD39aSL6Yz5c/AeVc5m0PWblOmjAc6EuIePzxnP/srU5qyxT+F2k+fN0
4mpYpgX+86xrrDpczY+j6QEhqzcoLMA+YpAMggnYAEn8lou/4+27jZDOc5ZsP43O
XQrEkctDFSozmy5hUo2lWyUH1c6qPYezyu7t766jkKQ0LZEZzSKw3X0yyMpNe53l
+6JW2WlUVV/chMEBiHFFyHMMegGwviMs6S76UGvcv66GQ8V9dzMSuSvzg5W11Q6R
IBtmFfh2lV5dtcSNwmvIjsfxRbBPYLUFx1Fxwn1NrZIvgTTGhe3wwYyOe18VyhhP
YpbL3CVSQJOQaoilikWaQ8m+aqSXRVJhGJImQL7o8bE5b4YNH4RURE4A5c5q3I91
rr6s6Ip8e//UJbPb3cC7AXOGW7nPad5wXJrC8Xg5Ufnf8oqieoM+Mte4DJFJ2ZN/
gtofP117ZJ7hP7yZCRlXxT6ErZyWtlsrRT1I9/p67uAI33rFTKgidIb9/s7YyrIF
ys/9uG7U8tJhUup5sRIDnkE/6vG05uJHm54JocaQ0E0ma+2EGM/BSNiTavuCOhMD
/NC6K5DfA1Np3canKlxkqQbVlO6YIjCFr8mW0DKIT27IBhzwtuYIBJrjWy9pkSeu
TWO7pSnJ1ZfD5TdTGOk9M+L08Lh8Rq9B0nTeG50Qi2oSlcvFxKQoOfdX7pJfyCz1
Sl6gO1w4YzrO013709+YYSCnCiqWKkmdibDrw9rgWDbmXigHoylzIeKvtqPF8L5b
sfsWgS20B9yKT0QqEbqfi9moub1DTXAcvealRhKNSAb0mmNDY7XkkmF68MXqP/Wz
E0/Ri4CEde2E+vfNLd2C8URP0gN3AMXlw1vzAL/1y0Drr4Z7lCXDEB6ftMEUDBFB
w9lvmRmh5xoO6JtuzHSDObNIC4NdZULLRPzD4wMzV4O/oPIr7aq2mdJfbHbHsdjq
QP6gRaAfUF/y6/71BnacORMuNgppp99E6b2LvnpoRi46Ax6Hk2/m7Sg0nBk96TkN
HX0oc1Nr81U/Cp6IwxtZEpkTWocD3JsHzsZCNPtiupolHsW0XXjt+Qc5tYjFrnxf
gSlWCPZA2TmXzIEOOYKlgXXIpPPZcxdzGylCPY6gUdoTQkvGTDCC7DbKOdvOWDku
WKqxonGOwSwHv5Ge31DP1o3jJCzMMRXvsohYk1/o27FuBfreP+WbHvyKr1Amw5jz
MPJLkIHMzaVxtsCLXjR9QR4057n8qrcDL7Ubd1+ZO41UPnawuS6IV8ABv1bkEipv
6Rw2Zvz5iq79xwfwcIHSLgz/AfdhdDdW6+5IHn4aviO9v+1oCKI1T8IrN1Ffce1y
Q21YHvO7OWTLFboPglJW1/IIS6OY+bQJaPWzp3muUNFD0Rh1NCa8fgvCfdIQivid
usLKCCzU2ngZPjOkf0TTaOfYYSq3ML8w39muliyw8Zrn8tpjRDgNuHyhVKmVoxnN
l4ujbSF84AQ3jwbR0iH3GX4PIag6aiWhzpKFylWGHHxBNPQPAOjsra8hDJjOAPdM
0vABWXYVWN0kmb/k1TwI1dQZr42X/IUDEZ8SAv0JfrLoBHuGGA8xDd3pDrlz6ZVu
POSfbxevyIwwgGqq1rgrq2TSlLGT6Ed7LMmM6c8kZQKoOVgWNWqE4r/dtCURfJ2L
lPn2W/NFn03za3phq2v2oG56jTkmGPOSIDfODK6z37tdtn2G/CI1pesXHIDsw9wg
oitJ7okxrOI6qCtqCOh7ARJgThxEJ88KAUWqPEKO8vV+EN6p8CWTFoaY/qu6B31/
4tmuNoluhrm0EDd7XpTVlz9A+OJ9Q1V7r1wRZw1J8jiOTVL2iPb/FjvLAKgnh7kn
x34KW/D1exHrfJ5vG9qqfKPrpaC6OwS3/qYQ3ioVjWP2apDY3cUl9BJJme/9yTwg
M3X5NPMqXBynLLDNi5x4pXOJPr8uhpdVod9X/zwj/e9BFDjuuZIKOhuoXPJ2n15f
xTTOw+x/LiUUigvpXwDRPMvViWKMNGA/i1eG7eg5AsYCewEfb1fdVp/MZ/rw1TT0
KXsnX2qaglxQyd2EHzZPdcpbB+pUAf/jmO9NgEezMy34hw6qD4mH7iMOoTFhOYxq
4YcNKcgbuvCDpSUlRbVgXFhvACr5/6M+VzM6R4UhvahneBfHYpPNozWiTvBVlYVw
eai3njVKaXWSAgiJFgD6Sfn9VfpEaYKyQy9/0pDlWvdx/G3HRozFRq0QZ5e3zbo4
dRxrgLKeLwCHZ03qcWyCbXrgxUNcUETXpvpo/4XRN65N1hYOk6KkmC6+gCV3JT16
48lAnoYicuke7c/f+5XwzWCkyLE29U+dVohW90PqaP6rY80k26mbIB+Rcwm8pIcy
aTI2jNbyAC8vFEInOs1gmZkw7atb4jVywGP0RnfLoQ1s6G3IY9gaG1iv77mhn6yf
bKN0o3vpjNIZkYKhtZRqD88khuZQR7MIrrsE+2PuTb9WBJb9SWySjV5Gk9nyqjkw
GVs9e6TOAkSrHgvEM3zI0Sb46fGGu0JbolML3/l1P/SAdpt36iTFNKAMPjoIFEBm
3l+RkpSWR87a0yHMRsPVkcxB5zqWPldCiLDZKr/ePWz9+O5xeDMixKobvgMFQGMY
AFweddXECdbPrFYbDKiJ95596+L2mVkM8WYvMbtz5X+d0AulW6TQHbtM5F4PQG6b
y0CsgTkd03kM6KFsN+2LB90tEgTgUgTjyzaUY8CbCV4MUVNl7rTdSeTSaRaDJgHV
SMD+aEP4KuAeAUbUfz/Uhk5oXXNuVmMgYZIMOQpFRgmkhh2CHQfcHD6EQ8ARR9Dj
W3XelXvBHuNME0hiQLrniqHYoIv9F3rXXbl7V88dekNzxdnjniuUusVN1PV9SaO4
3yjapsYTeg87CtNgcN5AEamU8E22CXEEsz6VjtHoy3lziCQDe3y4M70ij2yN8JXj
mJkdDD46uFEe8D9sIgxo6NJnsqTL16aUiI26x0IBwUbRfO7Pt2NAnm8n5ZhRchpa
gmP86Iha5K3csLyz9edmDFggW8r7Ir7atelOFIo1pa6FxaJO7mUaylG157BHaBjl
Yz8VaBYXk5UAWHxWWj4YCOCmS4rteogMOJSaRHo6qEHJt/Kxmpy7r/3QaR6aqpdc
z+tn7ef8vLUMmDYKHCCW3JcroGc+/4zWaAkvm+RgwoLRviVyNpwuqfvgCOtRedlU
zqCAQJIly0HifcuKDgx21LfRT9PiuZNSQmOZfsRJks28zFtm9l2ZYFmMShp/lpg8
lOsftSG7yTMsF7Z1a22fxzSgb1LZi2WCdWmVyTbGDUbU4UI+DMVM7uz13RRg+Bs5
gUzhvgMJ7gozBgvbvJjA4fz1qoEld6OGNoDa0OCF/QStNqiFdMwcMuio+GQYaYPk
5JVJDz0U19XngUQcklBAvVWZbV1LGrym+hlqCuUCco0xwaO/3awMH09sUxpzG4JU
TSXcfBXMxE3YK+KhDFbjj/siNTNhGe6jKylbJiv/kThXFM9YtI6xDU/yQdQG8xkF
iWSftzcnML4g+6Pmc8eXCEsT5UCoKnyyJ9cxD0adzbdcxduJg4BG7UL2LVOSlpGs
O4jYUw0S0yzPrsPxxDK+qHwjKcHmcut2zqb5bfkKnL74YMMRt0HjI79j5GELivtW
daSTJ/e3Ar9LCaRqVJQOYzSrWyHXVUBKeMFndc3psmOKzoUEeZJjAPpOX1rlBf1T
FB5d7Jdkhj4mm/wV9DLNL4QgCDowjQPr+XR5Mf3frn/TkFNoUVLtGRYAvV5uWaJL
qQ+fAxavJq8AUP3qfYsRSOlpgHkrKTFaL+Qq9SfjlDaURGd0nVXPeVQrGqQSG3rO
tUUoJgca11qsbsvJk7tCcCNbtUN2XSV2HpEvVg9NtaJ7uIbFx3sIfASCvy2lgtqf
7dn7VCiZ0STVGmLwnpFPE51zsjQw0w1jDNnZzOU0UQ41ajtoUFJfjeb8xvltsceh
W0+wAGWmL6BeXWZocmlg0lrFqbN697M0Sy1wL02kxFntkFFRyN3tI//1qa789VAW
49o+K3o5tIV/wygL56/6YngFtRT7di2l17OtNcpIKUnYM4rdW5WEab6qlGXu+bgn
x/4VaASrHaKm2sWxLNlkNm5tvn69GOFOnb38rtY5qLOUhpFzfAVVT96t4mckOxVr
cucJipOPrg8NKy3qD1NRhWzT4UILmEAWOfStK0MtHmf7GMUJMpKjq/axrKljZh5R
wDa/QkHKsJW3la3InnsRoJA785wpQgJVcR0EJTYf5lWQdwS8kM1Q0tuGK/nbPsPG
Qamc705ERjeVpVH57FnOpKh9f4i247fg6uf3CSzc0myJVp2K8Dh0ebDeMIaJD2ae
eKw+jtp7TxTpQizE45BUCv30AvxVFeZn+gvCAUkZgYxotTE11aorvx5Y22O++k7l
Jv3jmlvzT7RzIVRu5Flig+J9eyl63uHihaaCQTcKmOleLjuadSaxP/dlp2dVLUAR
9CXQ4G9a2i0iw/kFbdbowVSFTgjbTZyaJ9pcxaN+92S52kKlNBNYJ6tJhNk4seVh
At/fnVAIAluGxcPBaZeDZb9bYyrugHs7aDR0+gzRUcdmvJIBIbPZeNU9zI3H0JSX
ibregv9rXTTulyx6Hj8QQ5XXbOe6wBFirETKPaL6MwaRokzROpG+9acU+i9BGDh0
2EBiTuQh9dEQXgxRKn8LsdmYVuwtIpx071++yuedoG4h7OTjxwQrxqyH0KKaKekM
m+kpsWyA+AXlxV1RjLufYB4bZT6vdwC+c5qR7KMumS2/BOTpPk4MUWuSRkXcOb5S
Woc1+MpsFaNZA8B7EXqnst6D2uej6x5d46hhnpelt5FWfwbZWouoJF+y1iky7/PL
bTBHWBYT3k2Q0PYHBrGU9Aei6f3MebReql2fueap4ykP79O0QMyvnjuGvgAM+6PE
rXVa5RM1BmLMNipnn/jaX6LVLyvlOH2FvCQa2KZZMcLlLi5CInN0Wx26UZ3dpR/X
1YAFJPLfONokmb2SIWEFqVhBHqUbl67aQeFAskHczBhpEivmycJh64uCi7XuOqLh
oTcKXeftN2+zR+okD7+9U933hlti+eB2g1TdcS6HjdJ0+MFYX0uiqeb95GtObZ8m
t8pQ0F58GW0ckdk6A/BgmM6YExvm2qf+crpfKaI1IirnoMLAeyRWJh3ua7pGmtel
jMXrK7bQBiikhhVq8+qhSzn/csdAm664kn85JK2dyNPux8sHC81VvrnXZg8Xhox/
vd9f6SV3HMfPNK06k/0Z249MT0vHfk7W4pT3WPJaAUGPlCaNiHnCRReYxs2BrnUn
sXExTsCTXzqH/glYGPyGXw6PUVCu/M4ZQLpxWaz05+lCqqgznzFjLW9CBnyNENe0
vrAkPJr5leBOYeyrg8xbZI0k+u5yjKEdMoDwYMJLpEkKHeF365GRjqRoXU3LsByG
VbwZ2xEDU8R5U7JJudpZr2Z8bF3vRfoelA/pzXBjbty0Hk9xe16M4qjiqZvyGExe
YQVo6zBhrRlydQhF4ty3MrPc0sI1ZYDv7AdNSX5rrx83PEM8DLH0khLn4JLLGu5J
WXFWR5TGzo4JD+HmfZ8B97oR7Oacl51K4gIRfdZjZ8H1Rb37rhuFAf16J0YoLQpu
O2CwDRb6W82Jdw3XNrIJ0xGL8Xm7jh96rOWF8r8w1fX7uI6cxyBw9TvNIOw2wF8C
yhjlYrFjsmcKENWFIOcdKMbz4k0yMbW6Ql+RkzKVExzfT+VvoiBMRyWqnXrjsDAt
saWIMvDotoNeFef0WkiN48EveF9AZA7c9uXdBQKfR56TwjcbwJIjD/JfjC6Un3D4
1WwBrCcYIuyA9hQcSga18KS5lDdF+CqXghJD97UYgoDr9b7AMdZhvr2CcRdJCZHP
KtJODeYgeoVIGE9zCmIPMnqJOr6RF+3sVZaKhSV25XK1ZhEgmYV064VgTwEdq4So
lXmTn2fx8Bm50GbSwCwumtRdbeUzlITNNleXb+lnTEx5kqSazB5LJn8HgDLOQiMi
mQ1TfnBihnkVGNr7okb9vUXkiwtoBsqHQ45hx0EXlGnG0R2dzd4JeEaOzNkwf0HU
kbY6K1Fg3lgZgl9NhhKdQFCBdN0FFjp6Q//grGXRIMOb5ikaJHfAZC4lAj6ejxKC
bm5SFqqeCcutKYVczzsBX8jS1SQkO8Ab3w/uJz/1k6W95Ljqqu6aDVMFLz0gNg9W
AcRP8vnPYnEzsWZ4LwKE38/RMWoFDnh6uevqYGcrVxZB/UP2r7ggFWLx1eYjrRto
chzWVfKKo1tI8BWi+UbEelSmYZPtZeFyQqcznVhLheDMHmOuu9QJUKmnzjRE3SyY
zC5nJnVzIl9kgwNviCJlzpZu+R7nHU91Xiy4sxwf7Fy2KifxNKb3xltWSGURBLH5
eHpAnpC232vrxW1ZRZM4IrpoSZAUK59KLwYmUJsjJxph0lOfdzAoHWaWR19KKAOj
lVBfnBcqWJwtmEcJElFzEnq10D+oyfeSsTlGUlxKQY/8TnuL7AyKGGsVYjwxNIpt
sVZ0fFwud1yuHaCWRWeqchQ71XCHkAYHs5fvBNGOL+VYnboG3RiWfu6ln7ZFVf0S
rhxmCvcdNq/rUNLW1r2Z5na7JYLpSqbnmqCrFLrnSpgi+oov9rabikB2s7aHYIWc
wO4ZV9ADP6d+R34y0oR8Tj0TG+IGUXk1cxiDAkVdNu1SIXNahxIxamzAGNc3LJT1
jctmtVAJSXtsvt+v4ttSIYBc2/JVXQ53Ge0RrK9MXkWPHfZ8bkkMxm9pEjTvnRNx
ewJZuPFGHd/kGfGXscCTOVKS0RM+xfmxCf7bFhh2S2iX25JdtbzZ/KCt1DOayqNV
ugtNWxrygvFPwaajlawlqD58Q6IIFa92LSM+XMsxjC6f6UdPi3k2gohcHvAMV87A
CU6h25c85HG2DSXeYom1bcZ2+ykAnOiyl/lJjtHd4V2ISJ03v9P3njICKXVu+K7I
nsx1VqL8xTJMtEXm++Lxpq+4jDKJYu47tCiD4AVuQKJLe9c3ytxmt/ezMWgLR9fj
2mTYWxL+oOBzyHXEgagoQo+wV7Dh/AzOjyMM6VLuplfXMiHNidlc54JjIarti1yP
6j3oddXAubJm8MwtXwqTnhIkJ8vGsu8CMZtiHziWGZuYirsiL2SjrZ6DSJmOVCxg
RxLKdmaBhaVklsKwz0E2ef6AZpibtKW70pp7rxmCXqNz8KCAQkqPWWhMnaeXb27j
qJO1cUQ+YoJNWsYiwG3ScAFyxkoatK2Yg21/xcajKUbl9aIYyUhKDRKHIoNEoqAS
xs/o4sqEH0W6vTc/bkBC9TmiU2ktjZc0rcWebRWXO1fY7uRAzErb3jhPeJTGPagm
yTMt/tL1fOOO48c39FxMFF8F/zCuVx+9LibvgZUPhBV6hl5bK0jEIbs46MQfRozB
oXjz6AQPXkzfvCd4+nlgAdeDxyQED+BopRuKPJdMjACk3GUmpvkoW4jxkWSu1iE1
RirxY+8H+HjLvuF9vorZMG25AegbTJVHGdPCH1WxrQ7qnvlFBIOmG3psLiEkgZ2A
O3hal5BuO7OKjoxsZFPpNndRIpmnYGxEDqPR45PxCkyJ2Xq+42ooyanncQeIRhMB
HvyAU7Yp5i19bCr/BeAbI4TkGarA7UoYGq16XQNf4Lq+ATNzOcKHK9R8GUdfUF40
aQ7DxuBx7Wy7ZyZkRRTlmyBUA4FE1nQVEBh9zGlARHsgm1W4ufYL79Da8ixYRJ6x
GEzsvMqkfyfJgsjGb+G6AIOPPyWVQ86jzOmPIY8s5NxX9dS2LHKgKwB60F3DUSyo
1lelDcHVia1GGiiexz8e7INQftHSh2GYVHKZ6XIXPcChxacfVNPNe457wozlQZyK
i++oRlhzQMIufRap74uij6gmyE3T/lj/dVjQ3PrlzfguHnQdUGU/3WSlTfd4M2JD
5eNjdEraF9gLf9qcNBaGZWM9v8TYrYtEXWvQRP5pyipNUZMqcQQJpp2VogYY7sAc
PNL8S6jmYojmSOBrC/RotmQmEw37bZHSqrCJUigUSCuikS2l3mD39QhU+BCaV3yN
wkyN3l7OmIPIw/xIcYrJ5AjCvzR5lAEY4a/UYoViRS0mkZQWnlfr3lhlMTZ22Zhy
2pwDk7JKtXSUWVyXeju7zIRxu7chS2MPEBRn0PCqz2ZmmCgHH8vIYTdseGDtrHEs
ictB5ieunJByBJfo79ZSCT0xchomBzr6In1HfvrWxRRZDuJG7aAq6nCU767Y6rN5
WrJJW3KnWBz9HaZj0Bn9SF/g5OZe7BfkgHpucKsSo90vk3lGnmlvbGsG4h1RL/d1
5BOQn2uNecJ0Y6glqGowOYyRPFf3sC3ZIGbgpUhVaxufcoJU8jZhigY4vTA5Z7mV
DZmxw3oa9SM85bQcPZqwLKo6pCryVaDcPKjlJzD5g/AJTZvgqGludAzcdETZT11F
gKyZnErMG8bahOoGBUCdqsPE1GDLR1QlTwRESYZlz6n4b4QaUt/hy7FIrk/u87nH
gTVkLZ8OpySHkr1xdVShau8JMhNDtcM/ggprPBlI8zYigwEOLRLiHeFccbdeH7Dp
fGDkv/RpEPteLO3TLXPHuISY/bSOjd1peir/i0K+o/lXagGFrXD62uBxb09DPJu2
Q1sUlBxurBADpI5z+DTBZT7cZUuJcTVJjp6eU2hwL8y9T+Hm3iUYUFh47yodKbJc
h/qxzQb+1nu+bf7YkxJarA9SIvL7NJe2L7irg0ukgB4L802L6ypFztDILoC2T1iJ
aBkVULZt3Bov+guQv/Qgo/CiOdRvpcxxotj6uHEJYSP6k2P9ciZT0uRBBJ6585g5
mWciBGHenf7wh7wt1sGzaQ2SEwQDqlgkejAvRgMqa1oCOXh3maXazR7dvrt6wmTI
h/qNiBxDAEuVysFZlgqzwmViTo43tAo2V/nVaJm4x1fFUfPrXAT+RP4/o5UMZUgl
9M0pHOqrzKjHKc7ExwKLpYgV4BM4lfcR3PeHBMpMULicq0pdKCmlVxmqA0JUfzan
oyhfMxLzJ3Mxj9bb2OsnVuGiB1SZRhEfMTkiBhgluJ8qiOrMx/1g9IJ79mPacDrz
DZxYV364GHjhdaHOe8+54hVOj1bg5u+Eb6hnTTmGISSWNYfIWvDS1upvr5FfA9Nd
MKgdybbppN4Pbq4bnXcC9rGbvLAynr4jmNhAzSnQab8K8Ndk9KbZnCoW9XwQWh+X
JrSVb+NAlww8BIPffrl1HEgJj1iUfIjBnL3xtQpv21S7G4jLo6eXm3d8XNxsXarP
foobizx3HgXKP1pfNI8lSRVybywbgt89395dW5ZuNPaE+39103cUm5y5hYR5ucpK
dSpRB0mW4p4iOPrxMWI8yhuNEVpzHbm705tuoY6INJpTkx7L7/ikgv6+I0e8XFLY
xXmHx0/JvrDfjd4p4vqCi5WqDQBsaTksmf+nEp1qZay5kQhf69gvdhT8WWbcFAdd
pDOjIOs/N8tpdwcMCa2lxKHVyj19ggTA9E7xlNFL7D7ycB/SbyW7NtHn2qOZm0ji
LpCUn0HK+EUW4lSexGpTpUzVgLFpggVNGe702c2MwFaIrALS+TBuN3GKhq9T95vt
Yo63ef/JjNgbRmbcGeYQZgfskHiJDzwkCOEu5AS8bnyBqYM/qir5xjsM22mEVZZk
fKYKV3AYTTkJPa/s6EYAh+lSeqV5iK2qIn6Ii4YojNPHeuJOClcPxnv26Ndz+9c2
QdP/pS2zq/AGZ7GPLE+IFmuJYd2ObJg75q1sN8C3W5yCFdtqqdHn4f5G9zo/kk+V
HHqGPY+K0lXOAPhuYmaNzcBy8LQrxxSXHeMBOqNVyObGGLssvlAXZZodyRgNvqKJ
+l1m6B6sw1f4eSSE7Yf+oyxS3E4w+xHVm+EGJo2f4g6FI2mI9mgcDvzBScFiqWcV
L1iO2biyyTctkGs7o2bzoKTlqzSzwi1Prfg7T8B9V8TWRU6+WrrdYQVpkQb6Hs7u
t1HFFkcLXxeqWyNiHTOepvuUQiwCe+UEtRqR2XNXcM9ySn9LkpUoVVvJJ2Xuhrp5
4fEVqNgHpUaUWw5w7UabZMJ2WfmryrmM7/jyPkZy6D+1D1rvaLYCXiZSwjzrN/Xw
ca1s3rzbH43FzEnFnjtypzDWT0GmEShRVZZvm+mAmbUTuv+hkdsx6cwJiMmks8JD
o/hb+fUilVfI+Eher6NTTW7Vf7/WpZzRpvpoqCm0/p/YPR4MWwDucK0fYGyz6A6H
agnsCdu7ZeMkMCojQeE8GASQ68DQEiwoXcT7UUGisGezCom4ebvEknxxib+i7V+O
R9/qrGf1RcfGLvXL8PyhAKzTdv/EEYXv0Xy6Xhc4exOBFrDYehSuf2ialozZr4BG
Kc3vV7kXgC5Gas/cNQaKE6vFmhkSm9iN277/RUJhGj2Ds//PwKzxIxhAlHmnVH4r
xSYxEgWtxRLtGfVhvx5cmSjX5koILAuTvBnfmeNu4vWUt256nl1+IZkLgr74YYKo
aeSNF+Z61tjlwxasZKXJuOfRMl6h5MUvWKNpaEQCOyh97WHsORDpH2CaS/IzcDEU
Auv8/3vx0/TwIYEzRtPI5W1utFjFlfOdGEZe1Wddjgw9g35E4hxJdjeRr6qbFdZO
tynFRWkX68iqpzb85tOwJW8o87ATqUF4RvZN3k9zL8DeFsX7JXMLrUF8pt7SGkGJ
8IE7Gltxxb/pHhERWHyiRDaNh7jIgYIWxeIULMLiboRGXdGAjcz8oDvpBgEI122L
/DNz2ldqyoMzAS133zWftManqPqAXVRMWcgxmMQ1w30Sj9iWIkVfIYYRyWeF0sct
tu9Ia7ulQ/jL5GCnzw3c4ULN0Zw/vsrvsSzMR9D1HG/W9c8jkxXgrl0qiu9ijHKK
OUgwCfcgch3VRhnXFLaLPdgLXsbDy1S8zppNo5PfDT8QWzqe06/flW+Azr9qkw+o
SL5qdY78H63V7vtt4HwFV7PQ+B/UIZks6b2nen55bx689v1M8SJe0PR5X3jpYfy4
g9g2GOTlrCIdEnJt5HhRWm0AuIBZmbQyiWVHQOEG/YGPPByh+k5Z+FJxUYo4Xwgp
okKKHW/b1QNT/oreI8vvZFnxzbH1NW6dRhm5hUrw/ShM/o5XUjw3rjMgNc1KcUBb
/HYuW5fDPFFjezOa/l5HupmD07stegEeokcru75g7GAD/U7vQP05YBcfpHIv9R8E
Fe/usvUiZI4Lc1zIgtT/0urpEf2Bv5T2BpeXl04K1xT9pRO9YVzyYRqQcMocVG/J
VW/DY1PTq3tdrVy4qiVqkg/KjOq+Ke0/3uEfrHDFAkK+cvdzBMXnoQHOZPA6++5O
Glu5hNNDAAyqwgfLYabGTBsVmZqhttAYairs5qj3AH6TugNsqAJt84JwIcCB1LQs
gFAarfPKNxdCvDr07CldqhYBtXH19IVbgIh5pkM0DoHTBSOw5THUO0ypL+Y1cb40
1CNOH7ekndSX/1f7XgL1LhI+jqCL1J835ECjswyRvUtHPQTEj4FVXiIT0elba4vn
FaJKHfMkfDs+WDxgF0sz88NZLEpb5x6c5/wy8FT3QBXLQLvAWn91bWybpfBrTlXT
mVSZ7D7dQEXTmDybfhmzmoEbw+loCh2qVKY26ZRpwGBNBCXI1A6J2pom+5UEsL99
Te/3/01h6BRKcIcgRjo7Vun0tABC9zZ7fcmIMODV2cN++DpK/DzcdWvfRjmX2b0F
8YK9oS+rgvvV2wn91AITm0KaepVK7CYUtuc8g3vNP8fdIrHOG8IzR17T5u/FezkP
3kncy4ZP6+bdLim/AEBXtBMYUeaNIMfPu+aO0dcscAUNFwj8ZRgsKDT6onfujnHQ
Ehm2c+PWJnPNXIgsCEgrvfcOqWssAZHaoX1eeXQv9BpBF9KeL/Ocf0mWJkHooJdO
f6csg6lMEWWOMTSY0S4uCOVudfnYTp6JcS/mcgF2BoJ6Q1vXcRh3LOzqupzAnyUa
P5zMQCn4zq7ShMg2VAn5MRPtcUaDGmaXLybVGVSFxiLdEzoX5oGSweSpD6aza2/M
oP1W5ujG/kBk7L60/BaVO7/FJnNwVuvuvm0uaQpuVhz9OFYD+IyEoabAlFL6cmYZ
/nGFlVGoKGpj295QcQa+9QhLPxqTHugxiUKnfaB07XEK8i0cyGlw5MLFwOjqyuH+
iAJ+nG5pEBkRssZixm2VjMWPF7UUbNQxxrGPoYyHXkTBzH/+lROybV0b80Sdnq7j
+1ns/VA0EnHiF4PQGg8O4QoRQoBiUKtyEkjn4Cms/vS3uLTHcYi+UbzA9wIkC32I
l+RrOKfZadAfaAede7xYHHzHh8U6gnUKlF5MDuUGzvEFD0vMOHkaIWlrtIX5YtKM
9Ib/ZJJYUuKv0VWtHNBoSYstCndYDZW+cREaa0P+6pfHTrce6ignjy1yXkXylq2s
gIuCJ/yMonFClxSHsEP2KjWRC3qTOq+GDPGr2nRqANpKneZeLcJWreedzvxGbeHn
LtQPVo71FAcAALAtJjrDmsj+TzYrnYWbb7QaCZXaISuqMc0T7G+5csqi1wYHraWJ
91/OvXAcm+Vig57nI7bZ+SVlEsyqguddJp3wGLkgEIAcnbQOQSg+5bTxImsiA2+X
TbFUcGyd5AptkWp1YbFeU0VYEgG1OqBn3/VD8v2/m2G90v0JEGNaUnpXVBogq9Ib
RdTqp/Xga9QTqjMCrfaoLfxe/p7oaFBGuVmrH7zlKNS4Bbwo4XFx75NaN3jXGGQ7
FWNjWsJyL8CrleC+N7qUe4H+1CpWiDA07Dj0UCL1WLwDorbXRuULZEk2o6+HALQ/
X01LsjKNqEr+SJz8xEZyy+4cXy/8hEk+4E/QWR4TOnwOqAKqbhGmPBj7hm1XxlOI
Yn7UPNZl9RejO61nFYk18RAWxOfGPyGZs4BC/kD+uPmENs2LA6VM8HXNUUPh6t9K
h2cAqgsAPt1YXdf72TNuqMim7Wy7wnKocnK4otfhnbsZF6RzpiKwbKf4sznjgICF
zT1mm2kIToonfve2u+ascicNxfjypNihI28KqDTl+kJeSGFCSe3vb6SrMW6ESC+A
f9/0+eB1mztNS/4GuSMQD4n9BmzT5nwwRvA6AOD30gOrwnC7aT7jgvoytIVFpY01
UlWAFyYcGWCbzm1brGAU2MURQHJVCoob2158r2pO4VmsOmHKg3vTF3SNc3l72Zz8
9w2vIKa+aJNnK43LH8ust4z1nf0gMElEaDOwzV+C5R8PwQfAJfKJne3/BSkalyLw
0NkSaCMRFZaIP1xheQPgZPBagcHHBFI7tYJgm9Dx3SjZ3AxOFGX/zbOGacZw2S7F
x6Oo8gnzWuw+6QYjLTpbSK7opzDurFz5sAc0u6BM6faU5TZiCgSja6BHsbwIGZ5c
LQaD8Gm4uiMsYuCBW+bQy9tmx8GberjzhtpR7wh0hsc629MJSP8Qiy8Qz1u+is1O
mQRVazkZnAxLqFVfCeytITBCgWJZpdIzP5fRGcVXYyokqR1EawnV81n/xmFmCXhv
Vzg4Hr9xOOgyCO1DCag8R/IvDgkxcalSYkOFoGnYi22if1iDQMeKPxcxmsO4oFye
Ql9uVxEo+oq/Ahtle3GgHhuuDXyWtD2yn7W0vtkY+oHvZfJPhwfpu6in0N+iKyK6
h3ZIJZ2ZkYNG5WQahnKQXsYT318Wj9As6Zypqq9nquaw7PqDTTCxPHk0n4aEl5rB
ggPmzmIuNBWy9ktVXY/O3l7n/WTVeOYQhOYqp4fFLCyQ/tyHRyxOWzdfIT4y7vHP
s3nZYj1yYIOjSIovb+gfykDKXXPXUD7DX3/n5Qo7/l0O9YrUXMpyX1HY50D7iLAv
AZvlFFek+2G/gxDpNxHNYjl/VB7xAbguQAbCmXgHNzsqH/6d/I/HVGKBR9jJ6I61
I2Umn1UUuQdI9ThVxiZEkL+pwY9yR9l72NEAnHZMH9RoKUqizkOaTqnUuW31XuAY
sOy6Qv7fG9XlaRQ+NzNz5aInI48EjSA+AfjUeGfPw62j4/k5tIcOP0v89YrSHPpT
OA7dTpN0r2wZUcwukXAQNZNqG+0rFkKAck11GI4t07vY1sdzlwon88jTFlQWfYmS
9QyAJUWw1nPlU/dBq3bhnmCmvs7oTdtKKDTlpVKCQaiBy8MyazNO2rpUee3sb7HR
LHJry9xCZHdo6pIxF0cF4bUL0YdphKbGewZOtU+hWq/BGATEJOIc2D4x8Wbt2x8W
GAM6dXRFzdQ1Tpyxlu9ye5t18gIh5XFslXHCeUqCespqnCnhKgalpAIG2Rp7CuSJ
kk+5GauRiDWGIa8ZcyVIvWZfvz46NSPpoOpphD1OUiROT+ABmJZfZzlKBLSW6Owr
H6YiNUgmlHMZkqieuRssmxirDbRTTBad7+lqdEm/PHML8TyLjZ9W6jDA3Aoc2/VD
jD3I95XYtpuKLOTsjhqMx7fln0qb5oGc7xYRlVh5HMANuZhdKIb4O7JdJUjEJBPd
JJqoEnGsMSxTDybdPTPnTnElDEz2EC9gfDFcdNWjrcXzb40rk48OA7SraKTntOV4
voGTQH59tc+QHQNRl59KXpJNEEIgRcrrTJgypwR0A0fLgYfFzm9a3zqE/83IWDSH
f2tiZgcN07USe14bS6BvIEAXaN3bUwOKL5YM+Go7gYilpmZsibRkphl2jB9tNhi5
yYlAiopjK7GY2oqu74Gui6D6gnw7VVwC8oyDiN1k3Lgjqxaaxz1R+pqBXZuh9sjJ
PrYz8iim4wpILLCfnxHY+mZw9Ht4WRLzAl09hp7jeRCM+eUzCqTRw15cIXNyrZ92
E5sdpJxYXw/u1rRA8swdfZR1zx3iE86FjOoadiU0aJchJxMaUPY8y3T+RX359ewG
gAnwlohHcYTLNtMTf9KDpbjjgOOP4yIys76tIjEuim56Y1U4IOtyXBKelHDMi+WH
c9wln+s+fbcLt6hYNklvP/+2l5GYdhNgYPYCpY2fZK1aBL9URWi3zstO9M4iJFZQ
SSvTLAJoGPiat40FWFuj2QgaupCFCErl3UlRyE9+qXLs04Kl4TiqhkZCuuAEtpvX
CYIGAGdk3aX0AArtUYPk2J0gyX6stvRaQSr8Gk0iawyfdtNwDqFxNz4mTJfD+wnz
6e1mgp/xNog5F5zVCRNy0gjtFJoBmhTmkrhciKZ/rCdq47g+eAfb3gZ2lTCboByz
scRLW3JUtvx3mWwS2opSX8e6+51o4/oe4kJetbV6nLR72CALqSC0+rXPLQucGRu0
9KjeijDwIl6N2Eu6iYGQnnW3iT/u/F7Opp6mIptgDQU76nAmr+VTQXICB/E0/yjw
X/PDVTnc3gu5+nFAE0WoIiD1EFYZw/Z4TB7PfT37qI3LkFexptjTUkQ+u2j8yKMf
kV5YYreKCQBC37cakJ/W0y9XzZ2eYJYBLokrj++MEGcHk5ER8L8705DCoHkboJem
FqTaJUQv/dDQerjIlu06PGTAjTw5biPTkn0r/eCT5nQh6rFtcrai0GMMkXTMrk8D
d791usB13ydAQQHQlycOC8XMgmWVQwcOevV7MBnPuo2YSaZgbh0FhutW6hwUV4Si
3ZAD0VioSWk7+Ez48JXn3nfg7rlpyjQ6+k1uXks/Tgl34Zf586S8vYgiU2nNlO8a
t2S9/m46deSducyaCZ8J9WiY9LRxwNYhvDwyWFt12SsUl3Q+V16lrU+6wO2om/6O
roMgVyB9gG563s+N/bT4+N+pXZQPMjpbu7rzlz2Dewb75r6kgqVwG9hWN7jRszto
ZeZmvT0hZpPEZL/xPJjU3FDwgP8roZZSVtJ6NXcjegKQLmiS3zh/59f1MclyB7jO
SlX1qRBtfpXbP+zddGpnB7N2NwMpAbYH8JbH6RmAwcdImL8HtEAU5WmLiWhSrC36
4pu8edGCF0JW1lYDqv2Qivzt8moElDK4SRCebpqlyr4w98oHWDQXz+IPYE8x7q7z
3Nllusf8cgjyai+iUgIh069RO0yQinxdeldIvIMfv/yGSD99KFi+J50ZNahHo+bv
uPrLJwY2Ovr0Dfv+Z+LSo5awKxGJr5kTLjxHjHn3P3S8xNqLZLu24CZ3eIEVAmqG
Q19vnJxlyMLh08Sw48e6ktCk8XrutMA2nuS8D1WFEWHbIcOrwtcDrcvY0xU7dRUj
ggL5XOrBR7Lkkp1aUcBGux2G7XtpP17dT8IlJMLkEUk7yXms/MWEyCECG4S8dAl5
rIgw5oOOM+Daoy0rGUcrEWWGM/u4spEqpucQ4VKMfAON7nNylbZPmB4Lbzdy8qDY
GSIM2b6Ns93DojJ9GJHJfEN9ddMQTMOWz7zuizsXDYaUkkrBYm9+eBVLxyhop8Qc
4AaZv/6clKDgU7T9BjV5LaQ/7xsvWpcBbyRJac9Uf8p754e3qPCx2NzfcMeZHNcT
GB5G3Fle50uVZ1oZkCkg3LondWeBnWoCihsyL2n+KIUf4zr1D6Oy5Oic1ARCCXns
zZxTOX84JrdbNChIgV6wrD3z+mWBSz4fGO30i6/ukY9JZRHthPEYQVYT4UOp7Znu
3Fg29SzutBp+wlUjLYhHEWsR98whD7pKkX6irazhuhH6LPUzLkXnl5ezMMKJWkWE
BZtq4EAt51Z5DVF1pUEa9IB+13gmq3U7d+fk+QoGOTTDPPupeJbKpW/AolB/W5Zo
4Id4LYg+Lz0eg2lZE/964E2cudCmXNr+ISwNgEWCgUmhSn/tVPz6OmfEolKmT4iO
MtX1LMKzoWUEyPhOIPZV59lVZZzyps/ZjyXh3ZNMFbHq9+zXuRmvqUA0XAIs+SvF
We86/xHYTsQd38mwjymNmATPfCDx7ztVho+LIdahjGoXQxvNjEUSSf6g2X/VEDGI
++SxSbfYkJYY4QKqkj1WUYvjMeenHOLHMrKr4uaJU5xnEUq3BFsVI4cSxd5lfJp7
P9KFACYEa8B33DpzcpagR7mVbyGfFGJCF9vAZEfMwQa9Zd5EzL81cQvbby3Dsudz
JWpbLuXrfVG43lEIaodiByG+FSTchxtEaOHgsFDZei9YumGJ7e4w6FtULzwKMN2O
wwOWm3v/KzkoGtyChfEFVu0rODIl+Z8DO9aOEVzGdlKu5wzuNu0lv7MkKZVja0PT
m+1W7QX6265qXggBD7xUNONaAt6luHN3XrCKbX+KEBKOZAeA1+gwHt51yl1ETFr/
6drtNX7FrzkiuBjD5fEiGIu+pOB6Hgy0Oy2sDlf5MqdMg7EO4O5IsD9FhkDnpr62
An3dvXCiheM1pKsZr3PR953y2l5G1k7rg1FyN0nlzt7IH9GFsVhXY6aFoOBh7gVF
bqjz2hbw4fjz5HYOq3Em8qxty/FPxt6lqb0fG2tqReJTtJTxe++R629+Aad+Z28K
+M+q7AWEQN/D2Wm8Gj0D0JNEf1r3MrOxun4d19qeoMQAwtht4fb3DkC26h99Buob
8jL0+zh7hq57juNZYY5QJS7GHqagADzH7BNxnwjo2mXl2B+ryECsprBhOeEo6aw9
e4axG+83hE6127B63S/ubj7RcijYypzUdqhp8Q9ujba+MhyvUDYYDdRaItoZc/V1
ZN6QA1Uxg24v5EYuB45yYSsOqkz/eHCb/gHnE6uPhx6ljdP0ddkDyQLeHi+dhh1u
su4ENzG7fki6iBf96ervkXPqM0h69iaa2Owd1QN8tMqv24z90UbFt74DHiKG+f1G
q9ns3DaTWGxHr1+fxqGHb9k2jFqTIASdITh3YUoq6/ZK5mT6IvwDKUBMMqz5MkGP
CrFO2d0Y5CF0964nSRmlQXMhCTzqT7/tFRiv1olHyPjRxLYJtGnOIvcVajRZXDgR
1coBZgYhMccezze6aUOwTO8Vu9pMlEpxgANnYKTDgWwZCTzYq9mJrtgTfXmuhCWN
nA1Q9Kdvg5suJuO8AVKm4lIppWU5nC1KLAPmCYHCauXeYMct2aZDld/MjibcRUm2
pB0pDa7DYjKqnwvvhoxamo127FvxaNqP3BLRLHcTLzRQaODD61cuBP6Okje54UWx
kPJhU3k3N2qHDUqYLFhrJXSbE+289X4nGBaIHZgFzRzpgTP8ABVH9frgU5FVgoqM
mofnTBd8giB6JOAXGUEEfWcB+94D76+yQiTNAJVpzqz8rQAiziMuVU0K1lAQeK5m
zt1mOmeGDNSUiA+vzNkVUm3kYDctD70YCXCxLGP1kpH8FIxX6ZinjvIn9hHSPv1w
4GGsnTbo/riQbJFinoWaH46RBhDrSvWglaNRvLGnJh3P/pZ5r7/HCKxM4vq/cIjn
Dj2iCoT+aXMGfvY9aXAefbXQChh+9avxN3EqHjgLw3uD9lxLEcqjUkvhOFFxLCXq
TCOTy7jZ5rDoQZZbmrPqR3YPDhE78JWUGwFD89+Ok1u8lb8PW3geKUHo5xb3GMIX
+wim8QksLGOs9mrXIOjSqDAnfjnUjibcLUcwAzVJvJseu3wgcdIQp06bU0uFYECc
cWIoYhJbUSpRr9Kc6MxDVwneLkAZ+XG2kVSiflTY/jyoh7Eb3moth2+nJqOg5AWZ
dr/WvdvglwmhpdVfIdPehiUW/EbpLBoJVjzqee1bArL9DDsv51dba2YS9BJ73tpy
UDjs8LjOoDAGzqDMrYb/UqwKZD7eBx8Sv27bt4w3Fd/67BOcxz+bMco3z/z9q2KB
61j1GqpVmiU0NqHm378EvVHbDeune4vteWQAsuZLIakJRTKMnrmvA3KKMHtlkVsK
2eFxRPTQz2bU/NTwiBzzURsbudL8y0idMcCnyVHG0uqHc292ljms3BFxdIC04iAO
V29nIfeBEUlH6sUP5ZH8fJpQuy5PQp2x2Rz53zyHGqszKQhG7lScu5QFhlUyrjs3
hK7pVIy6wvpCYfG+rN3PixauljdW0LTnlJYdNZ2LdaZ8TBDIw6EjjnPuTrJIEtZH
NMPezCel5tUoSsrj19Q02a28d6/GvDZrl8dmGGoXxxmt0fJ14ZZzUq52msaYP6oX
y/aTqi1N8Cfr7aMqB7xAFDTzI/vsHK9qjZMqxsR2Shs851hoDg6gfyPM+JV5z37W
+k0BAHT/Idlpt7+6aqiYS42XyZ1CwxgYjv/HvZnQZ+n2wxUl9veR0FsMTI4VZS+/
lfZbi7iUyxILBPIiKFeAp9xlBww2vqlbNys9ahAoLZU+NoTBKsT2FuASE5Imh8Mo
hSfu/+5uHVIwIdoFboqu5pO2+bzFIfc06aCS2e9FaCBkHhJWF7IKn40OlLOmX4uC
bnPfartYFBOwpXNk0WZW4mLZqaf+Q0w1T4pLJJiaHWdutnB4OyB+hbiNE6p9eEXl
lO2FuaBJze0GjLlTKS23yCPO6sTFklrJFKPHhOBHfv8MLfXJGqeEwJhJPy0/odNn
l3eyUlJv64YzdHgBI7kXHhwmJx6KWUBVRnVraYKeqfpcFpx6fWRiTLlLHlOvMScU
44qFekXOovYxInIeeXzbIxrauOZeiRzgooezwKJEEQIb2fok9b5gAmmI4mHvxvA2
26eersUKG6GjW5zikpMDxfVvrCVtuU+9KUTCYXwdtK3SyenvIiw3CMo/p2xGEhEb
zsNk6XR1in1E/sBm50sg+wngYRc0I9l/6ic5BRWTgAkHNOuSPVwFZ2dW+knQRL+N
qAokDFR6pc+0PseTWJ6eST/QaMFYIktpFpu+wBwoWw6fHU/Vfep73uL4UvNdwrVj
7UC4EtSZj9sG1Qw7kqHaJ5NGvTMnKzhumvXSXs2TdQku43/61NBo9M25VPOEqcTM
eX56cSNJIvB2xgZUfkY8m26NAlvFOUCSwD8sh8PWQ8aHXrrAmq69p54VRDfNPF/A
diGDaD1kIwAYyGvN7zPYXZBIlwEaoQi510betoofL9TjQxornjxQLyaOBMm3YW9t
iozpCJzIuuWjOYFSmXE9rKWG/gSWHvYQzPgI/5MZDeQEaTvKxW2ckqV03tLha448
76vjFFsgqktZWT+QfW7/yoN3dCfE67NPrsbkR9FkCC2bFwNt2tDTRGag+D3y5W8d
yHNwho1lpaDpnQvRMafgV51by8vTg6mb80WWkO8+cCen6g56ZImXMBuAdKQDi/hu
VfDkFDZuPu+ueX3AuShTMtXzVxaoTgIhqMc8yrPlipom7fQMaW0YuYVnVqHH83E5
L2CqBLjHyCZH2FUYqW3iEc4Oo+E7dKRcIddCrU6XpmxUe8gPwgHvQyRk3YWPEJI8
gXie6Zw1YcaEz7NnTbK0ZNDjLRl4wtqC/l3z71KjC/JiZsbfLz/YILzNWD208hAM
REMs2MBEh5lFgQWIbAQEtuYH3UyrCj3XKplAqLhED96RESXTwcB+AW608AnbvcJs
ht9D++2TyTvIho4sLubLj6PxXY0iUsHF0/AXtrFUApMpevSCHnPUP/Dz6SQaloBE
ZR+UvOWTT7xtjbtnRiDHGkyF+HRFcNeOLZlUXghuuOlgaI+MyWKr+TbhuVv/T8HD
a5HDfieQCFFmMrtZXnuo6q2v6MLnDNXmVR97BFSjyWJzs6JONs/c/rNRG/7LAjVN
ixJJQkYEgDIu3bENqt9whKnRFuI6FULaf/cwG0/98IpA8E1ONAvkvSTy//Yzjr6m
H1HZ4GAwi9diiSHaxBU3PvRvefhMGZf38xUby3B0/W6lT962tXjtW54eQZJX5hVY
dWC4px0P3OYZRxISRmCM/G4hY41YZYHCqSfXEs2FOqNp7fjIs5sYgkABam846Kss
CtKZdt+pfQ92xJDNjNfHbEPqtbVlx22ECpPR/sU5YtNv2JLiiBeLRe7buTksNOpq
IDo8o93WMxL3uhr52K0vgK1cP9J7jwEBphNceFFcIB+YB6VR8NB5cF7eB6PeyZGT
fYmTdC7pirxvsef7K8vbSJf1e8JJze+Pi6HVGV2OYdA/qQDHRCjjQbdYGtRK2Wsv
iJba0IPskdnd1/yUBYUcPFNyu9ZHj9matn9lEFzqdSJ1qLy96acTWRAi3rdR8GD8
7EnbnODZo27Y2RLh7f7LnlPYMXu3bRjNGcFp5Q2rffQPn8Dgcie1l/hCDslenN5V
Zo+FZD+FHvNGX5olutWc0W9+pdKIAI6RK5f1p5gbHdxWj662Q4DPPtSAKiJCWzOo
iUSmdsI7iuBKZv0gVMMvLKqO3r3AI3DAtUq7bxtrHA+Op9dDX8p8aXAShUOzMc6K
ozao4zQ0JolXDGkNjgztE7siH9WpttJeFoyBBWoUkaOCSO4w0Doc1ZpdDcvZUdTQ
rSyoN+OMF1lppJXMkKs8r/ST4YsfnrIhrb/EROhV+HYPDjN8QUyOEMmniXQwfN0s
QuFjtizQzjiagkXQuKiAvWmEznbhXflXD80awYrqtZoDOwLGUFXaiV9gU35WYQcW
zT+ENnXRA5338yMMifpDAtzf3MqvyySW8Vl//zMldpM4QgCAiYa+7gAmtEic4kUw
v+uhwk4eJvhkwBwONa2RN2YKkvnWx2ttcAA4eozNA4nB5BTtHU9c5ixrIWEErMqV
uPnmAvgDtXWDHB+mx3cQ/HzSTd2xtln16EbvOnrfvOzb6oF0yMTqKM+bN3HRcfKw
5v2QL8b4Pht7X2Bkd5wMkX3/xVBPIicvGhvdJcnhucvEyugkC6YQwBUZ02FZ/O94
UoBCzq1X8hgh1z3TbTH54i3lDkc8l3Rd36fvXmFRrzihjz1M/nuXJdpPGKN+mznk
PffcYWOfcrNue2KsgRRt7d2lsy9rQNcvgRn6PjSf/SFWfPJ+k8KNHeaMMgIIDyh+
sUBfKrtSUR8WZonSven9OLzIn2KSopfbS/X8ykDHX4sDdsvcQkTDOV2AxjEaGg5h
wOGzQj4NZZXW52RzTSdwfkABE9KDJzj9pRBiVAlY/9GSd5QBN2Z3qXpMFb21GxLO
SlRpwJwV8fL5vB7/zYWq1HyTC8cEa2A86qlIvQKtYAyG0X53zmz7itlh3uwzV9gQ
PxhYygeGwkiuFQByQ15joMPoUTMxN58jpY77rae+btyKkh5hN91tJEumlTh6ZPj4
+RxLyATguHUWsc5o10bO8E4cqntjNcQhsKsrTY+D+zMsbgFOybNFg2EYY8uEs8yt
zwABNBFFL9gh30kbpDIKgM0nkQEAESujJwzUsAdr9vnODfy2SHTYDUmpDzN6ufMG
vcBWhHdMjCtygl8ENMYuMszD0/IkWEwPONwcLIKGCDNi5e/fZkeXBtlHbQR66c7f
OT4crXyVDlrvKqqsSqKkDotpTn7DrGYLASiixfhtr/SXn6e+UG6cSz/W3OC9xdo2
M0DN4okL2R4+bWYJynKg9/3NxwH4b3mJsJZMIoGvE0jcgfEdnF/sxI2ia0y+VzAP
vsxV8o1Gtq7ipfb+9qEIbUaAeZtZ9gUg77CVaD4T8PdngrcZtWmKVlmhfmEa+vQi
d73eMEzwyyRwTD0kRfgTaXmI7qz0TAMlKAH7aJBnRsQja5ulw9rQOsDaBaamJlMl
K6i9y/73Jnq4EJVjVlsJoZ5OvE5nzSK3ptgWSGkNx3GdL1pyS3GCj0JmdmID35nD
KDC9mNcXo0LKkI16+tIOFOmKL992CHO1aAgvhBVJuB8cJCjfhyBQ2LD6kRnbIcsn
IsWV4c7TqxA7KJAymdh32mzmfMwLCJZqdkz+RCC1dyOC6HgMGDBrygodq3SXzs80
c6jZiiq/UNGsYIBPin/SaTYwITttBajZveY7z/pdfpG196QQJS793dsNa6jd2Ofv
A5Jg6/IHXvx1MDWGYz3TLcKwrv0rFQncQT/qimkJByJWyXw0xPPs3mm17zuNl64V
qqoEliZpYJREOsIhmyO1+qbXFFaQ1HfGlUJLkzEb3YK7fmIdKv2NN0TNqQAntmwO
8iWyZmxPeSzUmsNR86X2SrwvxdmBgUzrd6AW7hD1NopgPm4Iu2DJm8ogSlsB8+fK
Xgdcdalx34cQk6cuVxukEXnPl2/cT4zODKIbXaDzPlj02h6aYQ5vm7/xwoSsjaz4
bb6+nLlVxMsbEm4142/By/l+PGeo5dYwp1t0YFJm7pyWKmJ8aog9NBO+gkXDS/k8
RS1Dge+dWnocDrx28IMJ09QEglmt253RnO0gbNflOgW0OywykRL9Wc8OWFk8tyUe
efBz/TcGc1NsWinAYNPUDTlDEDU23+dudFWgHcqWKCaL55U4libAWqUhorWlYqGz
MeCeem1t2FRn3Y1Z9HOP7rns9xyMVPdHxb1CZKQb6eM/jvZRywMdH2EHu5hLNxWW
fZKwbEsKwPLqxlH3T0Cc1KFJuJEYNYTtkFk/ZEQShcZdAAVuj+Ik9CLt5AKL0m7M
H1ILw2mQSZ6kfp314vL4KnqV7E41HENX6f70Gw5/txQM3e0HItn0TNceqJLfxiMl
D2xdLDHBTXM7jevv6mBSABrji9hxlU2DodGiLCIwzGxDc2jPrpYnrqNJW/0nfz46
pG+X6g6hYxWXcmlDf5vUn8GLaz6g/iXMotMCyJQlQFrXMtwXbI/if7yB4zDebGBp
JlBwFrW3miVcOV9P+w2041+Kg96CptTB029353ltGA5Ly5Z6hTESqZZYF0A/2EYs
Yv4nsh8DhKB8IodrqJjHkO2HjdezAQHhaQRhi8XOdnXJKOKXWWZruq4PbZvVL2km
Y9EQFa/g88/iVHNTb6BjMYzvdILRtgmGLqW8GtOLd9UtTwnuzTNaucjcJZVVCHSY
W6tNG+LAKwjsdR1o33UqOpD6ifD/RuMcKhBc2dvB9JV/8Mo20ftBcXVbHfpjQs9T
nvboC2MoxNxQJyYIJKW/MYCMplWzrK1I9V0BkUU3R+/0JPj6jtg0XJi28qfksBmh
yglI7m7vZejNoQYErGzYn0SLzoO3JOagnmT4BEfyLGwNqNcZp3FeFqhqrJWkrBPX
a3lZD2nTSUQ9TCPbpotU7vlmZNgZ4BEWhGJmy7Y65Dr/Z+GZzVUzZ8/wOgsY+2Ai
q85B6ACk6jZlQFiL3ta0GA/8NFUGqkdetg24a5qSmKIswf4R4z/U8L+wb00cEQmB
QiZFrlqGEWe0lTbvOZFXXf1AShPLmC30VSkdj35HoFBXd3pBTQp1q53wfh4GgIiT
V+MUc9umMORXTZ7v17DPQwKEGcjCWmN/jdU4RoLpxPUXJOdkUThkiZo0kF6vtPQH
yJJf4808ngm1bQaY4PwRm5ByVUsT8yGY1sbkB0h+F+Jm9eP31uQ9X/+vEazxkS6+
p8Vwf2QBmDGSOv9t1AKRIs7kLWihReKBVJ31aFUDR7MTNOaLnlaobqfX+mcPbw9T
GtZGtrdpmVUVdI5xVmliHt9XMdWMMPGcqcefyReMa24YFuOLGFTjPf0S3uF5xn6d
4oaH/aKjk7kyup2E4nFlyhua9EpDYbG8nmUXezhHSW+8uVBHccFOL9mrLayvvoUl
K6jKHcBySEstIL8LnY4d0jzRlD/9KwMBZtmNmO9GrwsFUg2Sj9kZESZJG37c7N0H
t4C82hrbZ9SFrBYk2PiTywztrWeAS41cJh4UJv+t7MgYFnlQH5V9PNQ6gVysAJOx
sR/gm78A3pR84tTjYHvcRCBzpn4lXCVMJYZJ0dtRJvo4YPd1l5Qx+ZLBUIo8Fss+
hoSufB4YumqcicCqPjWGXuhsOULT45x/GL06AYhfE998vz7dExjRvBIr6XUCnEr5
lYMs/RMmRZbZEVPL5lkMNd/KHvQj3U2GZFDYNHTGT3NKBwvsVgeWoMOo9Hd9kqFV
z4j+LS51DtLpgYT8Iys8q7iEyOKc6fNtnp/iTpgURmXaOIBFfLoNr4ErFIYr9GaS
cQ3GZgSb4unJYOkMiotzkbc62GwFrYFAvLehZW9zDA4JqHOWrRt7coSZv06zGBS8
wEPiKPW/8cj17gjEffEFJwAqlu2cOMHeq1/8sjrBXKedN0m/Ep9l3vqnAiuIVVCI
FAf2kqgf7DiH2T4advNTOKyTqWzUP/ZAIbTr2Muu1IBAr+U3vxRp3GJfEY3Yc7sb
/7AsU26OBIj9isj1NSXDOC1vc3+tT/7EKGc66W1+H0H7LqkQalq1mYBDc2ZD0g88
dJKgEhXViZ4XR85ZdcQBtrDT9Wjr9PoN+JPNFLpHhpr8QdlheU8GfRFNFi6rGs9P
IymB4t6LYjryb1lb8AfwZt4+L/Ge7T3e8GfS8FG35/8sVUHanLxge+9MwZjZKqyP
SMznGGukA6mOd3Glrsl6ZkyB9dg6cY8kE2aQEqmuGmUnQRBpBFfuWDCj6uVpgrc8
LwNv1zk9v4vsmjwDjXwRMyFu7QhIdsUvLUWQEOSRScHIAHp1AhbL+EWvpkiCR91V
GLFgKsa/hQKXsJiYd9+U5rAPckNR/GS+ybwEXE0YRLGeDBe4HmGSIxxk+R5OwEy/
81KKKRsPoxaMEfzWWgoYemdlgTkm9C9rCGmQALyDP9u/u4ULg354U6hkM5ZDwdC+
GUfWDRCClmIwbnjKSpRFaqPC/Zpsx2ScRlYuJhUboSLmVa+GKfsYETyJtIL48u+E
vkCDp+gi2axWDV+j8iIRRRHUngwejBeAjVexQB2NYpQKfF3Zgp6Fi1wvIidmmjDm
HomJZP9HoXDijqkjCffMYcB3x6581saqoutRkN5hImZGxv8fz5at3wTEVgJ31xFN
nV5v/5nLD1vyzPN+m8Rw96q1mJVctYN5QESzdUrmqKnbS1W1K/yvaXcVqUlHZcvB
5bz4F3X2CtSn/sp25labR1Q5HSZg3wUofiSBptmUxH2StjA/WeEJFucCLXhrJ1cx
ojTyaDjdDBHywLdMCjd+DkgW+BToCkVymtYR5TRH1kPDhLGOChpik9EHv0wRddmw
dgkFfl+eaZZk7COH09+8KOkdGHoXAaTciWO6tjYd858uWLmi4bvbBJsnpX73aXS3
9iICmL+8eJ31UdlSrZ1PU6nQH8Gkqk5e2UybKItGSkIkDaS2lT8aAreF2WNmuGPk
3r+a97A+LED4U/JSikxRcVILW9ruQJkmyEknPSDuvcncTybLeOKxki5OkDlht0x7
Y7e+RmTl1s3gEVVH4wIOCufHIm/u86Px1z+LKACAH72cmF19KbrzmVdzKp7xiTIz
uOleeGu/ovGFayOd8suI1RDJ0aUcSzUcLpuJzb4Jo/dRplabjd7wEqYBWr8PQ+rx
hy20VfiUu8AGy8SHPUSj3Zi9zH7xgGmLRKjZlpUvtU7xB69bW7gNCWNJWEfwLlrK
oaGj+TZBlAyKNTJBdwrkKVH4zhgQoyAsGz8AGFRGUdIxTsbFkYm3hoC+vK0e2YPO
3kJyvAwQD6Ikc+7D5nnDTeujk4t6zIDn28LtqZMgak//aMj9yn+GvBsgPJCzgI34
lhVXGnvYcqnA1kfA7s8QRaZ10DBC5y2KbYOC6fHnO2Nixv4wc1rkQIVz8KmlpXSN
BGrYql3pICgE7YOZmWX3eQTaaIvzbMmu7eEQlZv6y01z5e/Yd4FgukRw1LcBKwbq
vWXaz906TGYB6/ClAHWGBPU/SQMCagd9QbLZXvpbsD2D38LLpSn1CsQeUid2Eny5
M7/aLmajS+iNBAYflytvxjf21RHlKCH8VeA9ljqcAKk3xkKTFXflMiBc/2i4A+4z
qL14QkLlZRTlDWEWwke++wO7cXJxsJtPc70dbqjiuvVPcFaOPEslD1Qo028AmZig
4slh7BxgMaXbZY/E1iGOonj2ENyFLHDjbFUMM9uQGuaV1lbHCjBUjHGPjEWCcY4i
iJSsYqr/ghCfNON5mXE9yMQHICGmg5Ho140D9jyyRs6BshjQ8tSYgiCUEIhqKcHL
UZ3nGvLmBCjBfbuDyRuYGCbHNEAFEJR/atrFXHstZDcO/u9Wuz1cnPdm4PVawZvz
bH6klMcNwWBRjN7oDijwk/9kQayDhsSFxn+WaIoVkX1Evt6xLpkb93zNlWPUne7Z
xctVLIn9k+p8AsZNiUlybsHUsAAJNsNwHH3guYuc8utBNs0NdT/qQqOxwC9TZD4o
VBaUWzbW88AOn/UsVbrVPCssUX+MGLBsq6CZJTuJ0cTJXDRe225Z/L41eStJQ4ZB
WyJX4JtJKd8ZmZkff/72GZJxSWEXDdcM3usH4gX5rZW02vvAWi2vp0ZfAbdHBras
EJnjUpAQVy/5pTcoeeVOr0dkgspjVIpo4S2ttEdJHxzSHiv9C5ZNtUnUmUNYPPYD
cFz15qHJmUBWBe17DvpdBeyku1NQzxeuAkoJ//aZWH84L9yqHFyqxL8H0XV99slB
YU4irzOsCS1w7d5XMUmSfcYBLQ+S9fEW7bbLB3MCWC7SoMh5cXEYzzvJ6MTdly1B
/Xlo/nMHct77gZLZquaK1HCc/fFIHa4ddVkJmze6uFio71UGNcem1zhJ3Hxy2Y6y
QSzChULbETyxue7GWboyAQT3XlwDKERQQ3cUuoMS4uq4AVf254L6nCN45KTzvXLY
uSU4/cjq9bXL6YH0kwq5+Sk8BvrRY1JDO9rMVplK1Y4LQrfpAvZBTsg6tjw5hQux
BeRYuNm3kz2nJKaIn5Doi5QTyQ1iz6Oi5CwV5YUIMFyc8W1IwGM6Qzxp89/ny1aE
zO/qFlyyZl4fzSbUaCOTjQFItZB72+jQB8sqf2g8rT7x5a7YZicEJ9LZs5QEnDWG
o5HMSjjPE9lvASR9kdmk1B7l17xqwYbdzPwE5A/W5uAOLAmXD+5zgQoxmK72H56j
BtRVVNz/YR8ugeQPxRRRM3RNu/3bN5DPoHDWgB/koeH/KLZLl2pMArNFxaLCDDxm
jnOhPXwwVEuWo0I/usAvAEKjJV+SuUrt9sTsaNNovyI4edu4qWxd7xDTUeZauT3O
aYeRqgDgvzqWRWPYZrRh1p+EK0DvtmSH8G+Ko1N7eHzIu1vTXq/R4X9hMuULYxdT
eWhl9lDmEzlKijIOwMnM8Bj7ZANEH++ajFZQT24opduERkmXq/1+dBKY4Ja5gLgf
oJ5TDLAUyI1KylbrkLGwecMJ4mOYPL/aX5LFSoB/Dv10lWhupSCEiaYClQ+ODZz0
cv+cHXy/5eVmtV5QfNJ2Doeubb6nH2+ioy3YACG2t9CCSxsQKUEVniICY0FssOCI
Q7GPSJC9UrjWUFy/iijtrPZfYkj+QiTE3xvjo1c5AQqp3UnZqQK2dQFXZNrEqsql
zDQTBmtRGJBVV2PWxMHr4iVGi4y8bD+xvH7mIHsSckw6KXftYir5YTnZTPOFBkyd
NVgoWADSehhoMZK7eNz0DoCdq+yhXSGj5eaZ8Ocxd/7bVS+Klm2GpU/wpRSoETwu
HIJ6t44yCnSL3SUJe6yM5LASjHVYVKtZ2Ar7EPJN4A5B2dRby0gtxOmLsXaVPyHv
Vx8sHQaIPX7wvze9VVHcv4YjHsrik77XE1cjmef4H9ccvTN8hyHO9mPVAR3cR+fL
5Im8+mOL1jEvnhey+8PvLfPUWc6MYsh/VGm9qjzhS0uO71/bWjJISMIGpYUDDnww
AEBQ+FHsz+3Z3XPdgjrDn4qR+ih8UVWDppNEuK2DA3fhlVACEmWre30LOWIJq2DE
AarALaDbnRqyFFX2w/GyAmvo6CFWMtdtX0I5u5U0DN2vRjXyhkNI8B2FaiqXTbMb
ljORNlu1lESr1mUysWO1DZtoLJrd+LuXJB/CJH2RAtnHt9a5s5yV26RNr3kPksQt
TzWUEqNBB3brVRHPLViQy7PWaNKBGN1+EmvvGsJTYovHFkhcwL2lN/l134RsMhGU
P28RX6jbz8JhL7yyr+TZFp7Hj8cdckRssPEQ5BXILkzqlZx7ykLQXrigx/hZeeYZ
h0bfoM1mf52VfB6nSqaBT35rVy152WPvYUoHt67obCmaabGK32EA1nCpboA7Wg5o
g8bR3++ZQ3iVL/AuCqmMs8bUOrtRSvIgXKwWa8vHegJcm84G9qJrKR2OVVtY90dM
81pU16KkYtoqiETHzF8Vf4ai5f4p43jxFvrJ8HzIOJp77PTvSTlziL97pPjmbgFQ
4y1I+HN8g1s7T+Vw2ci03CDBjZHRL8jOkJuxhMUoid0CS0HJZyqmk9OlLaJp0mkp
UkbPr+yFxEZIJCpMCvbbD9gl65jFOCrj0WM1x+DiTucIX6qY5fuIXYSgja0rtU5d
O5Ikn/WyhRsZZ0QhV556kymPiNeNn3y/cxBujnSDL+DvJrP4p1kjESACBU4d5mli
vs9/ZaRreLn6XvOUVG0iElmVe62MGD4tbiXbwf1KT9W02kh/6Bcjak1i5PgjExSi
4jgnjOk+2DbWOfvZn2kT6fo/DH9jawCs1OFoimr/orHIGkkgGN0wSzjFnP8Zh/Pc
i/bqRzJ5ScrgpKlEWDsrOgt1sXXJshGoOtciIt9D97IIq50XJyhaNHyQaiteaLu6
YDh+uFAg64eJcgIMq5c+UtTIDZc/VdCflTr74ji1iVh7qFU7Ggyv/F54nsXrZmTa
eYaRW3IDKVW8CPg5zK1wmjYuNrm7r03yc49eO6CrtcAP1wY+rf3/1IQWgJRS4EN7
D+hf/U1gQdqNxBkxeSpVHsj1o7vwgfVBYUXiapKnkT2jwpSyCzHr1L33alp1sbaI
9p8GfKZjnQ+Oy8356740JguvqSGZB7c6+fGEg2g9t5OjxoLrxaVsu+TlMBFz4aAK
z3FvxLe0pVA2TXj5eY45sAAPR0zEBHufUAvc5VYUIQI3roF4U25rXz1GhmngoWxP
QZavmhcVl2AblpxX+8Dl3R2xlH+0C+Fbfce6ZhLSw3C9dzFwJoYdm6uQ2aiQUL/6
izvjgqBwS3z6WWJh5mziHYl4MEIvd0KDlFGAKswtJkvkCBHN+Zw6uejSM7nj8lPi
bsP3pQfBvUisoA9R3lV+N0qI6I/ik+AT1WA2mmfwHBqRyE7tNHxoR09cUHFbgyZ9
zsowleR/aiZXfuQVrcmrTIvzr+C5RxFLLWJJQfqmlQC/9PKc6TeEDLkoJ+1Ya45B
ngkhKQ6wyjMY1T2yqHlBdsY9SM+Q1ywvMJGMlKmUui3ErJ90ZnrsJtqgoV6DDc3r
NPHePQ8MBih87JVRjhbQTyZ4+40mraY8Xyo4CdgBggGrZBXCAeQhV8FB7X+UxutT
CrTR7/D37Ncj4qjEwFvGq4kPtiKX5PrlukhGLP17lhWw9U081UmBuhsh0GezBFaG
ssFEUouODJk+dmKcUr9+7LmXl2WYRIvZPTQprLZu9VenpuaWHKPXm3ofHQ8XroDM
lPAFmnNHbp7b++Z7ysoluXmLLTMVEWsH+bnASIqwVPx9s9sluj4fNdMTruj51UWc
VG5uGIwSeEaNULDaAbUGoQMKLt8i1skK9rolTw1fLdkJYba3FzyNH/bVDxx41vHU
4vhKpnSPWlZ4owzXJbEbXbLeV/ctr10u1To9WOUuV674Q31aDSKExt9/CPgGq8bf
TJTxvk1NZBsg75WFtt/EpuQjtMs/4LcX31tg+YmMopIgshQczoeq9OtmcVAxEoec
M+iW1ANH1IIbNW+TSvYipamyNg3RirFzrV+Hx70A3mLVhp57R4Eq6OPuz9fO7hoc
w/ovrN2fMu33ks351b76WHZgk6lUIPqAZL55SRjOJIbqX605WS4SdTTcsPbPWStA
O8Ldh+wCvlXAZIj1ywZWsO9xARO0wzWXQOK83lffm103clHKt36VeQPIKHbHM+t3
jS51E4yOJlcO1b62sOU9P1Qg9d9fIugNgGssEjoX3eLQmxWS5ry12yzAsnNZ7mUC
X9Oq45f5UtQ2VLrX3I/4r0EpaD9BE5NEwRbdqnUNn/XcmUPt6/uLkif81alD11Ec
1TO/lfS4GTHsEpOKuszbn3gRngaj0eM10dnODACFYf+mQncU6yw83CbY/PJH6V0d
9L6VaG5UrEmP22G8s7rRCKN5H6wr9ZVNxV+cHVL7wdoXrWjBK0+cleTHs3/nCKL2
JXLi4vDm4pwUJ61J/NQaBZ4z33ByAe8weKMEoHa0fRgVAC9CZjzhh2yaswKsBTFm
53pXwPhfu9qkVHCLozO2cdmJ21uQmbtb7axdoxjuWzb1qyVegNf3FPIVohRGuOMB
XjwSXk7k6RFSgbD16koA6UQDnTv2aSa/yJCV4BDSdgD1JflmhB1U0PGuKMDvOoHJ
nn3EWP5XjSVUxsnmbi9k059FMe8Coez9XNNsuxgagIUMQsknSIawc1EYWFTc7iov
oPF+An9caCJ2UGvrWQ92HfnjOSIOzy0puHbBA+MB0ltF4hQLH1VwVD88CM0vZ1HC
a28UcZUK1xTPZEebQpU3u+0sXsraEyqU1SI4kSK/tI3/t9m3pRLKljRrUZxEuyHK
RsciJKGXV6c24Y1h5VFKtbots+LfvdI4vmgHw0C5PiYxBy7RhAJN3AWxumpYPlGx
X+be52U/GqYQjnMmXhX3t8jGvK0MSONCK6bTj6aNXOPm2GUhPISx+LXVPVo5MfYQ
IO9H9ya+tSmmfYFQHW6XwJ2QU6VwimF4EU4a3qEala8XPX27qi/RTzVbjKoBZWvb
FrlCcVrnHkPIq2jmlvxi31ODIZ6atlQiMghlYbPN6+WKaLV24GQOm/qmR4gM73Z/
23kxfpLEgZ7QXb+ibjgYepBxvg12akef/fpg2DHRm+18DJ4j3/8p836RZBk6L1Kv
mB3eBOaCFsB20i+MRL7djRsahSj//qSuVSbsWyblUdA1eOdWm779vN86apdO/yts
nIu8gG0kWqO9MtJdFx5pEokAVKNKR/ykSEnKnAscR7cJJY/iAGcwXkiNHXFSvoXD
r02z8n+On6YnhDmwyyJvyetfIr4fBgNoWmd9TGXWFvMAwFx1Fcn5RGaSJ31E1fRG
MfRohwzErCUQEP4Zxyg9FGvT674UZaDp7VQMzlh5zq7BHOxIGnvDHskX2Gqevj48
ByDw6DqFWut0AYFB6/X1/9B/SzBppked2gi9HyOi7F5Yej40VEKWSQXNiFLIgzUl
14sCp91gh1r96g8RQcbMrSKccHJW/E6AEYlwTlqxgD+okcSxkbro+oJ8DbGf+afl
vOiwB4IX2C6ZQBp+93eGT7eTp/FXFzMXjkWft8O/WHmgkUYzM3PNfGN3amkDW/Lc
85DB38fqNHq/4/zRHF8bVth/EIkfyvin7YNjYwigTn4GEJD6/m+dviEEJx4zhc/5
4IVAvMVKCKN+IBBGT244LfpHHezdVAmHuV84vEhZS5CWDN/+EPYiSXtQ+2fevw+f
PBmfoC2g34FnvChDSrywH9vLWx5hTZUcsp19rypsSLtNwZ+p7OXmv5sIaZDMECg9
CHftyw8Ue1CaSk74zcQYi98epcaBnxckL48SdnbAtTpYX3XrWpLwsi97S0Tc3kZf
xuJ/wPb85wTFxQezpIbCNrmFcDQpNMrcLG06kCXa+Q7F6+3DJjWp9B3kPegzz5oD
Ckau4TCGUgq4lOoGR2vTIQjlC7TUSEosL6nns01MqLLubouusS3XLKtiSQq2jWlK
zAzzWiZR1Uo0ZYOO5swo0arC0spXhkEx6l6/9kz/iArQ0pA9JotWD3e2xO2i8z11
rcpG+3leHLZDZAXtAV9N22RLIgd2PD1X+u1TONcqyel/jIMbTfFkqQmnQ+OhD6el
lvmjv4aIhMtVa8SYt9sSqbJ18Ad11xp0PVUab/EZ4uzFy+tPdchBXuJHAKQJ0dm4
dJgpjDSzjLT5iIZ+DZmpaoek5PrFBgSMIVmqdzEhwM/Sb+uWFUUv4YyXqV4PzOJo
2xzn/UGONJlKTubmC71W+1DUHHS+Fy1iDJWibQUizM1yct8z5amRqs6fAg2AjqQA
ue3uwtpVVyafs7eXavZ0KJOBNbLRs4x4GA3qI06kDHyzeW87kYXq0hNbjnbBSc4V
SlOjQ6wv9ibp9Rry3DGAJ3AbLsZXHcXu7bdi4GGW10PK+qz4yrGfpEh/0/cnkXzK
iWDRA81X0nGo9CaN5nTqv3oZ17o1FOnsKu5um/fD8UDQTU1ELwjoZlzGLU11QA/1
xIXPvV/+uZt6lSuWBSOCROIwHZTY6uKUKY1hJdzoP86uSwDcYOu6ScF12Rob0YVW
7b01VrH4lVP8yLKvl7yK9hdQD2b404HdjnjTfwx/1a0Nx5Nb/KXoxqUOKsHSPRHA
7Vdc7MLPeTzRxDcQN7+sP16YbpKSDhje0tfKXrTOTG34rJAn+417eJ/zm+K7X74i
XOh3xcleQW97uEEDw2uArv4DsROdgVAiSm5s/mZMhzigoL4lHJpNYGHD2WAD9d2L
td64Ap6dOp99PMbSD/2ISM3K8mzClBAs60rSv9y5GvHMpLjWqddXkzrxAky1JPvx
H7yEJNBpAPsQuGm9wZjmx49HPQ4Tk+KHKKTQ/5jlOWACh0toSrfkScg+s4NKtcOq
jXEVlXCNFkEyAt2bKiMsOaQMb6TCqRhzShqBz7FYVagGIUpdzN47cpGJsBk0FjQS
SqiUMi+7Vl6n7WDSeogaqbotSOYx8iYJr9rhxUesJYngXqBMwyX6QltQdInycbKJ
5TUgY8RNoRW+lUsVRxsp8a0GDJnRjIpMw395lw4iIl+d8yjvb+zMrYbZbMN2g8fs
HijVoDNQ3Eg3KiMCSyA6695iJGPBfpxdgHs/13Gm0r/rMCZsNT1kQvwXFphi1cJx
T7bC1ZK43gRWrx44ooEwll7yZhOJ8OhF3NB8cEBajiIMUku4amY3KhtufTpwEoM8
8QUtyTEqib35Oc5GJHpG+nd6ebRzMXKs8U1sEyitQ5dFbSQ+3l2mRjLUM6m+MJg+
nyOjDI4nCcvKPNIBdeCFk37qxbHnkmzo4AkynZdzaiz0nrm6DjSFhv1H3TD7vnOM
QBqcJcNiA9eJ+OZG/+hHBVfE3XCzx7G9R9uZhgdHG0Cz1P+NEszGyXYnkPMBVKZc
I66xPnCG2KlGJvC65SZdqj6OGcTphmlxVte+bS8ixqBwNWAkePaUoCEhBO2/D5PW
M11oGoi9ZyQIr7qslR+ikTi5f6cM5zzYxqYrJWU4BzcUs5wTFwxsyV/fO0DHCxyQ
H9AvAS3xv+mu4nNpUICySQLQLzq+cu5+B5VmeMmXV9oanORfvoK/S1Tnp+tTTfnk
cKlcQckpLspXMr7SO6fHNcZGc0GHk6oJSQs8kgS23KrwTeHc2yXcaaedWxK4yh/l
5jCmapQ5JfSELqRWFASOvdxkcrqOVmUdvMfwGzyGxYtFr3CFvKFXU5IL0iDZ2wX0
bKDInEI6g4f+NYKiECj/Pq0tz8AKUKXyoRr0qSkK3W1vJbAL19Uao7oGDV6QCV/5
OZCdkAMkS7GdZJlUTz+fHBycIG0ujcFdT/rsQpTrpwsnMEQfPbyR6HcG8ZPDGwK1
KWt2DO9CzGefTvd8XwBLhhrl/fJgRcTtWr4VUCfW3o2G+Fe/Rfd0c2+7Die9Egt9
bpBOPCJiRVC7KFbga1Ob2XhlfyYOjR4eX4b/WOr7e4IRZthNNTC5hgQqhEIXjcws
3o4gIw32qU0OtP+DMnoeSZfc/zTH+FWc/SIaJBXfH94HccGF9W37U91XI8l4Wtt8
OoiJC+QD5w4MmaQWd3+B7zy7utP8CszipX6Tompg1NV6PfAd9fXXPDVO3OWtVamJ
fHelbgg7owWyyNG+z3TbWr0RC/yn1azE8DdYCAqxEmlcO1sWp7GWdxMyJSOHQ9OZ
jxsFCvnmzP06Bw3vavG1nd0+TRzmc4LA2ZzTtDQ1H4wZN+gqaNlR4wXqRJeJwEQ+
Yz6q8s75/Ht8v1k3RYfz3NZEqC5EzhxyccJdEkCVnEIaKx5Sias+a3CRtn17vhGp
SMIHqg2ClA00h0oKMa7CfT+c7vIfkjmdWVmhaJ9EW25Fkp8M8LHGXsqTdDZiC21u
Eo5cR3yd/suzbzUZZEbTs1TmjbnXiFqUDdHkErqCE++PGSrifxe1fyYa7IDXQhNq
nGheRYma35+SuXw6c6soMGjS4cMhAysNuYZxuPM6+4qU7j5AYLRQeCjFYgDYasZn
dWjuDbQi74Fw7TJtKfpswRaQdytVmlxcVixNI6gW1IB1TnlIL6hW8CIb66TMeTRS
gL01EjMp8YgUB9DzoszQJkrN2U+NKStZRduDuDnatKAU167Gq6LNL6P+RC5TBC1d
TO9IGgNTN6f49A4g/darjgpmA0kGLN9lnJ4ZNwCP5CQ4uLm5yNVvgH+EytcJlLsH
eh1qy4qMmpb+C7yrqXKJwl2OpZA+607farNQEAwcoKytkKCEg4Kxd2l9TXI21ZPd
7/vK8DRHXNuEoEVZT8uGcOiId0JLc6va19HhgpbC0CbwJS/RSLj0muMa3J4VINFK
ha9M1rEiuOIdMYSR8QsaimR+1X27JBnO/hZvHs6sB9jtRzCAUI6im56EUXMc+NHX
bMnX01PqOJVx7ViPM91bJ9kPIv4AUPCD9t62z+3WzVbikkW8Y6n1i5drhPaAmTOM
4T7IOi2aHIK7Frs9CHPpegDnA0hd9mDXVZRvZMEiW7UKO7OxpewenHSAIuMBZnZ/
xkk6ASSv/JyXbnmta6BcXAuUJ03X6kw90QuAHA/EvgWoxtdfxdMr6jvxb0SPjap/
yzE3mWzfKV2XkHq+RpMq/HHxER3ukOi9hp4rQVy1xX8Gk2aFyXdZoXkZNwWKXW0c
9CfqM96RsxtRkNtdnDIKGpAG1e2kYZGCgeme0mrh9AiwuyUAvwEO76/rt2K2e5pY
0WpmNTyweLd9W+rZV7akTlZzifYfqEgeksPBrXHfveGqjcHajFu8lCsArwo4kks4
NyetFLBT5S4PLyAppO2Q7XgLLNsFpmKgFOKdgaXUCi7ms7HgyfmX49FRhvSLsPOU
l6QW1TbxuEOPKBiFupEEwGD1VX7MgOgtBU5O+8SQj/LlZgtkgqP2EmerAY4afZs/
TQ75gjoyjGYndCIH8A/lS1I3p/011rlhQ2Oz8LnwKsY/w0u4sxUYNadyZcmCUlws
HXK9p+Knoq4TH4y5QFPvSGD5VZvAU+Zz+A61U3fIz21bZ7pfF/aNHc8l1z2bvxcv
S/taP4BYT3caEH+7K7WALIDuPpAbpv6/JrntAPHW+dTH5qP72LD5FkPccuI5rEr6
U/zFLrJatll8dGyd/rADP1779aYH5o7iVVejJaxMv5pTNrlT1ReEUyiiLGXlA2Ym
V/P4wL7MVMCCkVPGxKhy9+dHJ7UW+WwoSpy7Y0NmBQbL28yUskDWk3KQc6s6/mwl
kqG7iwJG5kUq+ScGiFvWwiB7oyDszOo6bWI5lfT6aINGvGvpxaL/0E+iU9yUkH5R
KkRJPflyeZaKzlgVH7hrCTKo0jM6eytex+RUl1I6uUu5bfkVRzhKnZl+dkgGOqRs
chAP5U8/r8NIUQkTYzv55G1595J4wCrZQT5rGr+tlQJQHN50LfdbmsCR/Y4WA8+c
ujJvHoQSGm2W5XRqrR/Cj3AaeRmvymqJUeTaYhSmwK3gfoBaGC1+nAn1GZz9ynID
HTer7DD6S5x4zByBmRST9OlYXU+qwOxIqcmMd/zmv/xLVwKepFfN5RBvVExvzoEA
FkJNFyIuV0ce1b9Y56/3iXEJGPmKXHNV61CR6diSkhd47Yqvb4Qu58u/V5iWGPdT
U2WCgg48YcZO6wp/DgfNNYk407K+XV2dsW7U2QYMTh4amn7HYmA4Bkj+Hpb6Ona1
l1WAbBc+51P1qPMav7XtyRPwseM998vttgW+J25mzMu60kfdqFsVNvV6I+4/Pcyz
y9s634VI51L+AOOpSrgwZA+M/sUlpLsLwqrMA8+IXxlkbkH2nCHfdFRRNfwVvWph
KIqqnIzcfdErLZD0rpOka6xJmPRmzYzOIuoCrw9BYnTaQmJYaqIU6ahlBERZkwG2
cRcHbt+luNraWqGWFbUHP6cU5xBuIUEcLRHjnwoiYuCharB/xowF5jDAuXMjVW2Y
5bTqncT0v+WusR6Z3o0DUNzy5zos2/tHN+esn4sF7bVHUTZCw9kN+Mp0c1rvXAQE
w/li130SphccwAHYcbT/KBkLykSO2muj7+kH/l+/OnCorbgsDbMtFcI78Tq/X5/K
7IO0HsKyPp6O4wTzxvGd3z1tu+nfa80Sd09ICJVACqNQwAlb2f1lfqlkfXqFYEFF
o/dugN3VS75GcKYMako9h/O4vu2EbAyfgIMkNr8FQNSi4Fg6S4wF95l4XudRixyd
I3+YE/0yVfdrnyw/KRQbpFPVGE6wVxxYq1xXJt/4TaGUz9pS4ycJsZgmkE/u3B2h
cAxuZdW1Wz9pkdXuaxwwIp7bNHXFQCJK8FKexHk986agGE/hj8o1XZ8wUFFHQSz5
kv7s4y65Q5D89uvwh3N6vlz3StuNgghbSfDnjs9dHYExiEkrvd1l3RrmKf71T3S0
yb85l3sFNvXNCjYSsZdBe+sRIhnXVAPVZYJ+7w4/lt6Y44Jc9Rh/zQhQtD6jvBwe
pqc22dV1/S93TQQ0NKoyW8+A+3rcocEZvNWwlznJWlgNltgRCI/5jK787JE1fYkR
KneWmtl/8RWP0bAN2cvxwq8NJP62lITrqFG47ASwOggw7qwszYHz9GUrW9SFBEXQ
bVligcELEtN+2cSpSSwUfLsfZFPen3nPtDvg3AG0GyEwYWVSnekyMM8lgyr+BI88
kidrnkY7eiB9HDMXsfZOgJyMzfa9fdqSwYb5gPJ0gFsBiIuznQOR0xDA+GnhrqrL
9JSzwc5Fg4CxG78q2Q/5eLSgnVaikpmWKeOLbhRt5rsLloBf7b0WXL8n6wDUtU8I
GKTr017hJjYSoO86Ab5TkH4y/xBHDC3wdPoXQjs7ZxjsdneBvAEN4vSU6pZooUQ1
fNtuXnjUycP5hk1bRNXrVsmNyhDeWznqpLmsh0WrokMCjxjVBXkZcMPq1mjbWCYG
gAF8NZkrbjApWf2QMsaeBQLeB/xlUlpE8o5JvfDbS4jelJNYpqxGWPriMilUodu0
1GOVaN3T17f2bkuNKmrrTgGZvVMoNiByFeZWw7vrPXCSbeDAUL+PRYZeHg9jzUst
q+tFK91umolARUtADv8VSwJi/s8Z0rGg5w2MCK1qanDWQhzOgeKQf9QZYJeilsff
eoH4izfMIGlNigMiUs+d4Dbn0yLe11B3ww+pk9JiWMPoEFyhDqSAjQ7HrmEbqMuP
6xyRTs8kIxtfKPgaTHvYjkPyhZtQb7LkJVCJthIylPgJQIjWTxcK5mgMvKIWNRmD
BzMFJ86jDGMMms0d9uTvSqUsc5fEw+2tj8yApMcw/zzpBptrqmTsIIp/pzln5HJW
E9q1Gc38yx5RjuCJSpVu7YNy36ghB40AS3lwCaWGjDkyURIX7ZBlLvqd1qYeoXf9
JP8e37azp0ee3z/Zdv3nWHjNFLvjx9QcrET1vXFyn8licl6x2VoH2LPQafEYBMdh
8zkRLJVvd/6gKtk4d+8ug1DF7msjZmgHiHOmWl1vsK1DF9A+z6O6IX5BZlZZYUyY
XpW+sLHUrdrWXrABDLJO5bLUz6YyNpZzWiyIOIMcV3StDNpgB9Az3najUGPL5o2g
yku/xXe+rKaggFzvshYgfnvtAdUFt8IfqyJ7Ewxho/18soC3E+XVWZe9iMRotjBR
9GMjSyz1FaNIsU+qj8xJM2jwZ5bPFPwv0pZiuQq+wgi02f8MZYQrmfcIJi9eO6ke
h794t6LCu8DTaMMBNatzFvykeC5U3rmvZpGthvgkL7oFkdVFrcMWlsFT1vudlQ6B
2bhAowW31IklKecA/2/Htaf2thGYq0XN66ODaonmSjciy1wFV+QWItlWJAT6J8AC
dO/Le8VRp71Ifu6IaPdeHIHVc6HX2WUiiSbJhpHwm96fvOBd3kB5n1rmbdXvLCJY
wMRK9zT/iAxyT/tE6pNFG15hCWz6IdrhTpYp6bbsH7Qh1eI8DMNY3uLIRoheRQjc
Lj0f+ESr4Xd1vw+zHjTe3GV/kPzlnxI5sOMg2HNR2nJU6yHlza5NQMJJmEcYlQRE
pf1EL9qS7htrLWEgG6iZ8HGVCrJFgUpEmi7pLUR7ubCLkgHKb1DxpD2oVXcVqZNB
beG2OhdFt8NZ+Zn2NNTA6Clk3hPY2ZFk20QARQyR56Ma/EKnc6goU6CNQug9LmZi
ndw2nhwLMOfV9Gs+Wcog0ZrQC6Cy7czG66Tup/SXU72Ejz0nhkTpQ9ivoR3E+6h6
eggTrkj+um+NhPFbFeCFpN0s7RgjEC95WSg7g8GLfPfsGvtV65DVbcLXTF6SH8Z9
QgVJqCmUbSoQC6bcSOSL7ivSD1zctPNnCeVR1NQof911iNO7A3QxfLlaSoqfT3M/
l7XdVo6h9AaMdQgA8NcKr6DXz/aWRR45hzOY44MKAOe2WvCimDkJoPrxQ86+AbjC
7eLtwqagRLar5p8POLTue1joT1AlrjX6yOPXm7Zcto3rXfuX2zK9kOEMcbBbreJs
cVhp4wFwcovZWpgzh/eja+XCJmnH+IFCi9EYuU90mZc/mHJZm+AW0JNoOut7ID4J
/nQnU1dF3yFQuPtFKmgbI8K38SJIg8dSpsYAM41xpKDjd04jcy3pnXky/+sz2hfK
C1OazCVgkH+f0owqKr2dDLmXj4M1Z+3tG27MgAdbqQURu+4ni77+OENv8BcsK/Kq
MUeB/WNrmmksep3aQkkUKgJoHXPBmUaDZLSh3nsjlIQe+cPq+qKvE6zphEdUJcmq
w4jhU0voIjdmjDhJcsnqtlD8RtVKLZIlFN3MxKtFd91K6TluvgK8TiR+OJIPtjwv
YJyGvTaXkoMxcHh7qcNaFQ5KaF5tipNYk2MR6Hv6zLhxpJ5YaBhS2V8D6NN937jx
HqBXK5HdZz+DADRJQNsxlhMeXw7HA6muHOCyitaZQ+6cb4ijltyK24H1BNJyPajn
kHGFsy2d7hEa8pBJQWynqle3Aqmyemx5HN3jegw7aNxbJ2gj6Ro6+LCUe7MY5wm4
lIkpjqf+owXxo+upbW3NwRpWXOcGlb3cwhDQt25hcHtLUh+HTu0yRn0goNZys562
vmDN6DLqfXWa0s5ilhoayJaiLThLRbLaECLqwg/ef2Fba5FAFfMzB2yHACneENvH
8XVWrsKPpprPw1I3I2pyuwFD21vZrvmZc00DNq7UOzp2s3n/ppJr7p6YHDPpAGvS
5vqu94hpSTXOsKkrVf8BgOvBh+HhDHmxEtdcXomTFVSODyV0jxpchepILwTTTr+M
wB1q/dazVYuRAf5GTfRyW9Y1F66C+tGR6BVq9gF4ckNeOsV+VOwdtEtX/CIfTMhn
Qn2FMPZdfhff1niZQOt6ya4Y8wAin4inQ3RGh73VQkSUahSYokrlYpxYLon1+GA0
ZkR0g9y9DHn1bELuk8XfWqWesHz1vRO7Gm7IuOMzV4jWCu6bi6gS4l+yik3F1jeq
BYhoGXE/nb9fTrDEAI2UYcg/NJfh5DfhbCLNmci7spjkQCUInMiZEQiIqJeAiNS1
bI+a3NA5KP1m9ut/yzpEh82JF6KfFd1zpe+vsNGhItf0w0VS4RDjhwfh2PRe2SEy
VPHYiOXLYzo+W1bgX2rP1o3mWzBCU2aVmlJJNBJ6JTmZDHfpqD2R0hhrbg0gfl1r
k2ziI7LE01FyUI7XWKvWHKC8sEqEzgx0+TlUFVBzJfeibQrNox77Z0cl/7J7pIex
clu4AZO5U6PfffUc2BTpS1LMU/BeCE/c9Z0ruW4H8DsqgmW+uX18DeK0hvPWPZxz
fFXjI2k58iJXpOIbFmB1A/Je7hk9UhHCkjnv4e6TYuqf9ivtPF2Kn+JYIc4Gf8aa
4lDcWCsQ7LaKrY2GGc/egTB9sANE6iuJobjVq4J0fgyPPxsex2mCybC6x+zaz4u3
FuZ2assYhu4zA/1KcMmurUt2QTJXZcDJIlLlt9uYf/nZc3nN4vXdB2/Gg1Fiw2bm
M4AY9j31xdqWlfuFoW3ivOGdno83FFyWi7PgN11czojn/IrK6dUnyZtZH2o02xZw
itn7W6yDsA1bgxSBZic0Lz1FYnZ5CZfh2ywfTU+9G5oA1TbK/D9KYtbuu678gK3C
V3BEsyHRCjv6Ftp2VgV44ssOvJYxso+lEbh/ooqJWmdBX4G4fi1e34+EoURoaYuo
1dVjoS3YrfvtDF/eC7JKVz38jNERWEKqDDjp4UQtxwL1RPQ8kprExbCb3gQlEke/
BqrYcrPPQ4QUVMBm8IwJEBjRDTP0b6N4mMHnYsZEr4WRoZJnMcbsbJADjlxecEQ8
FPFiImsEwbA9235OTAoCIWkYAWYQ6aedIXBQqx2xxStqrrwfBfHR345C8eOAS6uw
t1M8IGScsTHKc757iuCV4gMeZZrMcLJPcW0A4+fpdqSV2UpnNu3uUKSINPGo0Igl
yUFnVD6APrwwxPOZJyYLLrZSfEmYHIf9NsvSTBLEY/OO/2RTc27fw4CMRhddmasm
KYOa9mth/gq/Y8tBFnrQdN3C27ONMx5QWaRnUr/Z92qZA967WJCpy9Evn6Teld2/
eanEIcj/QdB8LDQn9eaZjfNoqbHnVzjQp4RwCivOQvWKHTEm+R71uSY37U3VtfNn
46yMMzV2F2ZJzDseZgJMiQPJkJrbgnN0TCL6pAlWUFMgq8+HuL73B8UtKV7eQbhq
lTJLMLgYZAkSNcOv89HjnvTEyHjNj3Zh/yna8lg9QGBndo3KeLQoFsyILWNXwq3Y
HhD65d0A2IpKtx1mZbub/xB0XzD7GD5VJixac5xlD2aVmAs9UL4kkXXXrV3lb3Rw
gr7Fu2cnX1YHPtmUTr+iTT9SnIh5qQ3zNx5Ipeq4siueESjfnWzNoCLTGnJ6zOdn
UyCdp2pFF3nb1McrxRQnJwoo+5i6Uf5WOdeUwWwZuCxYyiXr+YbUj36ydM7hTXXe
h/KV8d10it++dci0W5sKnFEISVZt9W7UvXh0agCiziiJ5OHYIypYaRWEXBEv/7GK
0Jle+xUGjG6QxcvDsrqHwgRR82rnL6PG9s5hiXRuzL/WUHxfyUyYULP20RVBBcgX
5NgzhjCZb5yo4oZvJEnspPLIxYIWxeT3rHDjAJCFEXRYDdSdYBPVsxfw4WjU6Byw
YV0ZwLkVXzSe8WyI5eI2pNdU4pPGOCmocgEfBfFUD4LAhRQDtKBkwJvKfAZ7Kh31
aNynjArw1rd8SZowJu7KWyuywQIXH4K8/kgI4AVRvfFLOocHm3/KBaIOyKn/Hykq
icNrDaMryUTjHgqFxbt1gV7LjpC7EiRjQB1Aad+LkgE5NAaAk5jjKyt+OLWxEy+c
v0GsynaLAv/DkbnDfPo1cFH5TFpeFP/sl9WK7OulP6VD0rjVOMB5bf3r7efHcXZh
amjsVkDuSEMaSHfsCdX1t+vQI/3HoMSpAkHNWxs21yduXqy2PoFSCp7i2QmB1hiY
nld+9wYnu0BDyo1gedCjTnw5xdK4eh8CL/FiFLKstw9TY8v/I9PajOFk9ssdiZxA
3CR/gLMNVoyqSjnqqFPNx89h6kA6v3enHZWLHko2fdUcWbnv7N+tu805DBcBwCno
D/f8OUN8ZQVIWGqPhPXVC4JpNAdLlesx6DRVOmxUSxBalbfPeUN6nrCMbDWU/vM2
HOuN/qj7SO5MFvugGRCg6fOOLNQBxx7l/wW0lvIJxFEmSZ6+ludmdLYIHKy1d/5S
HwG/pVVn10CDVmI5Q0Jfy8j1bdsGBDWWB8Q0eam8J3366zNAb25mcbu84wxG4k2L
FFjb4Nh+y2CsGFx7U44nLSJqC+CjdcUOWK6x+ujhM+tscz41o539m9Qu6PNgI1lC
0Dz0LFHKIwtES+vQiufYoh17d3L7Pv07eKzTMPlpjGEyqd/ujtQmyACC3pUfRqur
AXeWgtEw8PLvF30uHMMj5gYlnZLnUbBW4okv+E2EjlLUhaPiiPyI+2YZByh0J8YJ
nWJufkShsppv1NH8UHwWBzLAfLCCY0W1Wn5QNYYJqoXfGto0SHby4wdKolzBhCCz
LFu1IDTuYi2Nxt6gdKwrKM1CxJX8z2dsKZH1fBOwB2dlI+RkDz0sByApPvWz2Z2/
HYfjT1Xgp8Kq9uDdP2UEfalcKwbZ5D+PYG4Knia4dizAKQlj8nkgrFfkK2FKDGBm
XlsNyXlWg/REd7HxgGVQ70JI3MZUxRDpC8KTR1IpYj5DmD4PxGCBH25R6avzlk50
PweMKCew/e83vBGFMiJ5r0059DyJQDjto4H/JewVI+ySAP/2MeF0ili6SwacDKec
IXbOR4nPh4uHVOwW0uCJB/S+4BpvnhGXwv2fMr45T92s1/3O1EKATS546d05CyMA
YEjFldlQIN2EGPa19kraHWJa4Mo9HRbq6i8YvKsUkg3SwWzaB9zVLK9eYg+yUCCM
NRHpj/UOkCxfOyJX2iOrTfyqH/vpna26vVGonbLtEoTXyspUC7Et03vhYmvgFpBD
NIm4SYMLUr7tTO3ZcTGrb+zCmF33KWWLRiwgpsj2zZYuAmW8PSFTB1mfeWqtber7
o6xqgaL5ksVZ1o2DXIJvPhhV4w8AI/dgYqtjBbBIXLyNIRwKae39JPcjLhUU63JC
4HXPBlhxFZ/BaBO9XbYZ4XgOyP7PP/ytpAApz56NyzkXHB8mAkzp7I9RS1QPZxm6
CLAz02gBjPD8nz99O120tVED4V+nQebAK5D1op+OPG9Qm+URyab8pum3/iZcVM8V
e6V/wVfPinZVBM08aTVfa58Wiv5lB0HlY8IuGvRTRp3HyJUgNA691tO8xWWoFH7s
UhuACE67MzOxwhAlnKYtk5urkoLuHBaUs+g/oqt+8OB8yQqZ2/K14C9bWRupVpMI
NTf45K5iQbW2k693VAWVvEu+ju1K+dcycHnPSJdik4IHx2cALs03GkCpDUxFB6UN
RIWzR5toshnMvlWQu0gFO/04CnaWbsYDgsSyrWRuw6QytmjX+HIbzphYGMWkPkwu
Z7z6QYdR5WpjlfrazVJbYgUIy7mjLFvN7kH4YP8ZJrWwfFSryr6Xu4VkE6kDPbOt
xGqilKRl2xeLEg1pzgSZq73Ok/78caQ81Cte5zGfhLEIW173qMS4f/VG03nP7KDV
066bh6e/GIpEphPRt2J3li8Glvf84HDN7xdMytUt5DQaR/oJodPtBDhlpRWWEI9T
vZA4wNe7mBONy0ZTlYsLpREpPkP3Otn8guWJC1Nge8VDmcep51CnfDGDxZLKW1N2
jn2uMcTT0CbiWbrP+FY5R0G/Jg9Ocqv0WlZwPUlAZ7WEEav/4AwWKxCFmvvRbkKF
jxHxpXQCoXjGT3hJOlrAWNBASDNHCBkYVvMdRxMBWCoo4m83bBJbMildT2ncEAh8
s/Cf54K0JpqBG6DeZxUuWbEQdhz4rl6viZvV3cvPdV16n7YN7K/rn+ZqEkqgJQJy
m26hOsNlxPWoAlKcQsK5ZH0s1xet2S54/QuS2Eu5/FScFfj8pJP18cbxLik0RnfW
tx64w6V06gnAQcqBINhmnvIPqXRJtvQXBz5uiReV/a5otu+aZYvsQSkRYMgosPAS
brKWyYMj+5BfRBd22QwoujC8dybVYP5JsItyQEoQkZIu/mwfzSYExGWpMWFQqcNL
wgRsxNhgvRHq4exw8bdbYqqhEcLHHCZCCBP8skFFpSXAaaxpfp7Yx6I1glgkYQzo
eX1sx9dJG1JU+venQ5XJTPefaETpxh5Cj5gqNK7t1vwFasxeRXOV2b8xRqPuNpHk
W9vyFCP/d5fS8BBRGlISAb5jCDZOxUP+EgpU7InB3ojLB/wwPPg7wU2QwX9upuIA
MJxvpMSfPe+02aol7D9anJj+P3BXgCXmcOqGDYZW+HjCQu1MiQjvAiC6EAIEOYls
r4zLHR1k138vBOY6Z57byJD+SnubDAeylFYzUAlc5EZOt4kQ80lGm/smixqcjTMd
X5ofGnWZySYijVFbMhtzZnNK0fav6TZH/QFCb8EiUuH60Agp2x+cqe3Nf+D2V5qu
J5elBbP3NP/8elJycoHFsIH+lyw/grJS19+LsrFH3LZSW+lByj9Djc8MRnDD/uAl
ViMrwQLlZZZhNs8Apd4ILWongGZHLS6TGFx+bOCZVH011PTulvfMs0u0D0rb9u9o
8VwSFeRDpV6Jd3GhAOqHtuPrhziQW8HmmdAtyzSSDGGuuUl9PoKf7S4noQtn7Vpn
xjRfdqCZzsJvTvCY7aVNQNdq32QKOGjcLY74HlUAVOgTC2EZ71mNSuCEtsoi1/0n
Q57GXP58hI7pVTmpLe+zmnRQXEmVD3B6njiSyiNzlAnDsHaJ0u9RojeM5v/DeC0f
ZHFK9fZGunZfuISihIKFfstyI7cdkXK7SGh88kp7kMdISH2KojoMvz5P6cOYFMw8
8mEo9Ps/Ahl/Ppl73D0FiCUNvJXgZP7aG2S+UWbRvZiJYz6ZmsWEa25Z52f2GhwM
dMAZk7zJiPzeWWtNzTj1hJuoAILjSc3z8v9bl6I7HYab8p0k8nq2X2BZmxDjUze3
9n7pBpDCAmoPJr7osm3cRb1Lwtng0ZLgW693HeOZfgLFYCxHIXr1hGNQeLVbDDF3
DglyNPjpm+9g3P/2+QnQ2nLULjnaDlpt0klkD9eQiMuT44upRZ2aZ52GgR6BViej
qOGJMyBjfHwlRpREOyVlTOZtecp6JSFbQe2Ujl0jtdYvcvemrPh6t6BJESfbFuH/
2nw0Ff6fiREcmsNQF933PimLD2PK6nopbqxT/g4dyZnrP+7KOoQF3QrmBV4L7QEd
wDAuF6bx8Tfmf5M/LMeBc8r5T5JnLc5270zRwjj0ESQRW1gU+mOhVZOhep3WvXA5
l05fGVOGLAhtBeG0q4q/AvUyXeUXvVYkfhTfJ+vg2Kb1ELjlJBkJmQ5uzJi1iFPZ
MFlfRW0cn3u2l1D9VC1HNABVWL1dUhIhTLRyNbaipKs6n6aMKx+HkpbhG5wNP8Rj
GJYBBDzSA8ZtwLGuSQQf25L1df61GRwOgMRf9w2pVfFRmmCAoc/HYPLjVBY8n6eG
SNp9mfQz5MCfrAUKN+7ymn+JyKRwpImthnOwv5JdmJkwmvPGudDWIHuOyusqEjp+
23vYqWnigU1oZl6FRXPnh7ZODaeeO0Kqp/Sh6t8Z/5mQfWBS/9ajt+psHkO4kDYJ
8Gg7iiuwsXMW9x7r5IiLZKRuVyt09t9ApJIXZzyBK3hSTyKMybhqdSCJvl/W/6/i
Avvmh2cBX7QWXxBTVeO9Ecl09VJJ5/g5mAG3EiKNoFfekB8FweN8J7F0IYeKZQqG
4t5+eJGJYsUGjmILM2EXdTS91ZcUEeK6jjqLmTvWkv11TQpca/xWRLni/4e+UAKq
QeYICjSFj5CQ67toXgC+prvkliktWSmbAX5dlpRCAkX+sdTwQJd3nhk6JYBOK9uE
wr3MLGYnyzKoNJF1lNfobVyCoTsHW/MUeKqddzE44H7Oavg5J3WVdF0QThqrdUBc
Dw8IGpjXZFOLBPSdu7KB6lCZWE/DWY1sPt5iR+pqlFi9Zl4gRWFnA1v/IboiSCYw
+PUCLdwh5j+i2jzxKsG/koLfewiIBZ5URPsFQ1776sGeRPCCBuzkOL9T3KeQ7l9J
cxitdVdOPdBUo+J1c8D+Z8I1IbkDjkUPJTZ4IM94820vKi7gMqXnXtJdjOGd5xxd
6pg8q47ixa7sCB7dOI/nc+TJOeoA0lXdy/QCrRBvxFop79IV14F+5G69aSxfvTji
fyNCaG6wpiYquuwTw8DzTZFUvRQxO6R6w6RgxrV7/v9sPE0WV4BJ8aXZYMXCxGcy
DD1eoxz7TGu//8TX6QlGtRQlFvgGYleAJKGRPEv2sbKFlZJsvA1xysWdZdeYkgYU
4c0JyH+SAQic0ykgdqPzj2cI1tu+51seVune+DEaHfGt43GYruWKjlD6qP2gFhOu
ihxP4kiZWR6ZR1hrki61PmmMx2YPQMXtUlWMdptGeWpTKohJEmvsSUCi1PisQQN0
OPiv8of55j/e3KQhPT8XEPrwMf6+jAlKssDZEFPktlLAqd6kevBQIRODDBZVI2aC
RNgyBiuTKdwfUq2Aoli6JPjBeWfwcfVHxhZ+ya4HZjNnfizahHssOo7kUXtCL4zK
UJ9BF4DxHF5gxjif7o2yNSAWvyu33Y9Gw585MoN7q+UOjVsEoelolmbe9c4pCUhX
b/l14Q6MVRIZF9I4MMQ6kFNkAmlRqOIBMdt3xRCp+seK/7XaXsxNwTfylmMiyf1u
5pcZE5ykRDiOS8uo/xHE6ijJ2UJxEU2dyIskOzVjo38QYsbJTL940V/bd7Brz9ie
Gb60Yd8XkI/BwBB740GdatwRgs7j05PiWtlmTCPftZeMUZkz7QTnH5+mcvVDABJd
XpEcS/O3WnljXDBNCfqCi4YXSor9WAHESKXaKWU0wOHpRU1YR7KcG47WPJ1OMqc6
LGaZMvOjZ0+F5xZRyYzIGAsDioNhqOqWUI8iTHeWdO3URoq8Pelfx8mxszh3jnBo
fWEIK2vknG04F5rPhOovmyKOMD5ydzufmW5HMsHGc1/kHN+cSI4HJudMI0WQq3rk
gNhAkFjqmnm2Xd6FtztsxuM6MtiC9WdmgOqzKa4kPzXwl1z8+qwtUOSZtRgL43nH
87/fP8f9OdhEr+BMiO/zr3My8oJ+Ov+b+pv/RhxykvnrjLNmE4nHPvXE7GnuoySj
eVE3ige+pdgrQ7dNMBWtfsXFG8XArB7WrPn64lzJkreoRyKzigkgDD22WzYYSU9b
8iaKeEk+miwUdyBFwuKnp9SQEf13aSxO2CPo12jpfpEE7ikRlE2NpufBGMijngsx
m8UoM1KZs+oSsFOxyee0FnUfHY1AI3S4YiUWGy/yeNTosftVoipJxdyNwekidOTp
DaXWbjT9AMMuqgkFeknmtxBQsOX741V0aFoA7X5I4EMNsqhDFaURODPBO3uIstKG
bQts6HRL54356ScAsjCvBcsCuA00YaILWe4XPqLgIMtdPvlkI8ylYXdFuAnTuKK7
Fyxs7Mjn/QDROBstCOb4c6Q/w2BdtfjUviGXMfyFCbDaMNzJpUtwyJrhgdwYp+yk
CoPdDZZb9MZabL6P6XgmuSu5nGKAlsTCs8JS32ZTxlVF2la9FtXvDtzLGHzLRQ4w
WQpAgeqTT46qNMFXQlhyXxRy2eI5WQn/zUULaeCgYFzXrGYmPPMCxgAEDAKeR0CR
R7alByMvZ/MutANJoU7g+tiiqtzo2y4OG0Ra92RBEmKygeUfYtRd5tBrC7wuhfAG
qopaTYET5Le4IH5Xlvgdjnkb9Nl7oc/Y00OpOLdCtqy7ozlvGzxeg+Phrhz2ifR8
8LL4Sko58HuiGE6hJXkpRZIpdOLfGVAG5IwcfJmDLD33YyXlRhNMghWnEeBMNMiq
D3lSqoRjdLgfAmvhLrowt1zzQzxhoGKooSe+STzg+2E6Ssxxx3Yfksn5/2K+7mZX
2fXHexnVykFH+AsE5oVOc4Vy6uLJizGc080WADqvIkHh8TfbKa9QeQdB2YBRzJg8
FQ5iqAUkbAFQOzuxIbZsOIru/uK++8kpONvVlBpqY1HcknlZrlYagiyJgoVEMGzB
1LQdjzKVBxNq52qwwoE/t5nOhw85M5s3vRLGnEl06fSQnCKaF7Oc3rgbh1Sw4pBK
TULCyeOgfDGZ3K2uzwzj5ATskCxpP4sP2cQ+lc10KrPKnWAreedwpWYWkvv+06bc
IBPSrk2V7EF4mQPhBWuXJntAU3S/tCNGvswTiBPuIofXOvnxadABLgZO6Oo6esfV
s1wvMkOqtJI4ED5XcU/G1Vr9pm6f1y/PBLHg7Pa4bWopFNJKx7mvim2+1KLLNeM9
zslxAzF1nyMRcND7f1Zyhv6S4j5zdAYLroyNkIiC+WY2gPRWUkyWmfrPsni+Sdtl
OcJ5na+eR5D3/qwI4X32vZzc5/11xe6Gp4WwoEkSrZkaMi9Lp8bSFPEQv9s+ZcXU
AWCORKdapOL98kO5WGY1Vp1Xpvr2nmNp8CRNHwZrgscSSjhAJ/yDGWA8v3cy4hAp
M10KlaY+6vLIkt/ge2oDn+eON0jNY2jMlFsmeFgTiRCq5eQzNEpaO5zodXPHYXoy
PBAa7uo1kKEfargJ3xB9h1XKYkbG3u0YlSEfXzATY+VX/mVMRLZ0ER51JUhUG+Xg
B8LEBxkl5HWFO28vBngKEDUU8fwx1L+Bnb/L51HBLqBWQ/bQCTDgYS3ryWIa9o9h
KyGBO5iXRas8q/lCQ1T5qvBwIYxbpR9wxPMpgwiAnUoGXp33MzEdIaCkmUPjaMS8
J/84/cmCuG29RJfftWuUMnJCvfUCEZTQahFXpnEndHDhc0J1rwxccGhTC3+W8vwT
H7g2pM6lkgTB4M+wApDsLLwoArPgRNnAmSBUrOaFVwU1vWXXqG7ELTCNDNyle6gy
Aj4mGZED6tQRsk9itc5apkAxXET2bn93udsX7az2IIvIYNR8N/CkSaj3n0FAvnYI
w6hXoNRYuCkniEbb/i0XTYgcG/4XAKmb2qrVWXYv5FC3brArCSdMzaGdynWZuPWt
WHseYgaaY03xKsU2tVnHhvhdGYxVLvQHeDP9FQJEdxBIzuJYZ5H6q6SMWhqbN7n0
Czu0IL1weVGJuVphNabmgukTRudVn/E2NP6UDlnGv3MBvb2izlSx7NfB/OQ7Q708
iNgGxsseaRsy4ziMnTMtavbXssNdgZZT4gAS/bhiKhht5uIpk0wb5ex9iK3PkP8N
EF1eVVVGwFC6Da2gZmMp8xPNZeBi+XrUyRnELQrz3GYZH/8+qj5hXlkZJy9Ftce+
rwOKiLDW3gMCz9VKKZY8hB6Vrnj7mIQEX/vTWgaTg+mrTV2EOWNDaHkge3YqzSKe
KQFn6V5gOGopZfxRGVg4VTCEReLdR+U/eHnNSfpt3vuOCCTbjobl4nZf3ZAK0bse
azkXfUhnCHeKPPkJMV7c9U5FaqalHMg65wAU82Rddja/yplHkZ4ROXC2aoYI80xR
xbDD+/+r7cSEObebfnk8oy/GpNORVkh24+TPFbg20W33lWy+uQl3FEIJJ9p5PRhe
GxGrKXMFUAXl8+xNqFmJglzOV1zKCplJHF8spxKGkOJKpPVAmp/O6BPRaDNVxuxx
s9aUWvY7gPNDlfOybz6VI8srgQQ7PX3+Z/A/IZaW8kzX4NzzD74vaa1XVEnMgVjz
CoxgcPI9PBduJZORxv/aJs05CDUHmdgoc0lAXoyGosg4r4DG2vJJQtHqZ/z0eJOP
T6dqgOxq+euriZNJcckhA5gmAQ1sSEohBdALCJqo051ZnFHNLuUGjQl8C83/8wwY
uRFVwXn41WFrBAoqqLuYbF499CL3XRiG9jkdw2zCzgsOFfg1AT37EQuRNG8B6KMS
4un8+U6NQG5xmkMcbSp32F8HU+EE2WSTWIGLaaJRqBkqBF7XsKKXlreaqT2N0Fdf
qb+hDLQ7s1Y0yXNiEo1a4FkKrXpYXcNzGQVTA0Hbcj6M+2yW/FJdzRO/N1JuCIuA
dVl4xTStsNOYjzqJsF3gONXaCPseBtH702bcBpaLcn2bQkR+9zANVWMagO89CAnN
OjDGte5ZXP7LXL4F1CP0KewuIDmDTQUH9c2ajTrjskhHQaGioEo0MMO7TrKLPGT0
HBw8woKPdH0oIcZhPEZad4LhysDKuFXpKzNz2e0MrixedhQCg3DkWrOO+AVF+kfX
2R9woVNnvoSXgSfkIhn7uVvFcbR1SJxySL8SDwgU1P5ST8oV0Sqn/qEPNgTl3gL3
aGB4Nj7+1tUBXH0SdLDN3XZ5dvl6SZz8o5V9tOo8dPU/TokDDdiHw+SJxoODLLTs
fDFyLwU7MOZyszc177nz+lZTzvUJQqfz0dUESb2UrMGoMfqdaxYKpckMpj0i4MHy
ixutMhPnfUfDh5o9Y1S2MLFeQZwwQPghJ+OvKMbH8w8PxtWguqQu/XlSwqqPVO4e
IGI/j8P2NuFW004L+8L7MkQ8jk5QbzqqQmChLW3rcchcovpDAxCa/5TJH5ektwid
hsv1ph5SmFJ6S9VLadOErcVrBetrihN3I2RPlrnXF3BUcth0DP1o2FpAdxvK1n7o
QIO7rpoz4SytLeNyEIkfnieOTWwjRlLvWFyd/3g9UlUpUZI0qYpBc9OzFflxBfEk
0wwWX/RAoRje/sQRcLnyOvgEEblLOcgG1tJoTkklFTb5bzVOgOZBmdtpWABvc0P6
JXIojlww6ZoHJ9Vm9beDF4joJdqfGFBCoHccL1ukC1nJkCDvq+JfWzokrgvw+9+n
j67F8wqVkN2z7KMWeFpaeRba7QAwZvjRY4/Qmcj11+u+eeF05hF/Nr18nyWpLagi
eOXY6lxw9/HjvMvyxIsvZr/aOlLwcvB1IR7/3tAlre+mZxmrd+WpLP0wVsrX5Nuc
xrJmAP/yyiJa1JeKQRWr5qpnDgy9IUjjsNL7OExZZu2URdJ8nWDNojf/hc/1ErJN
erIkg58juy5+D8wv+CALcEH5g4ikXZtw9AFPFa14MElcDyOSNWTALumKHqn1syi+
URCp+VMWGc5ZGyzxyDjEae21KuCgoFykUxgRrh/8bJ0/78+M3/c/qOsw9erOJEWx
3vf3+21SI/tUXXN4C6t56NfYPNbs8XMA67KZJvOVjdyBni5LkN7LnMSPaE+wUFN8
Dxl+p4VfnApLgV4+pJNCiEgxStSApl+KosWlrR0/D6QzOZlcsFA9JLDIXZYOwNpb
du8FtLsGnzcJ0QOy2wzKhMCXvPdbiuZcrRHQvroXOBO7YtiLX+Klyp5VYNsstgOn
OLXrl8/KntTwLSkJ4GiHhzjObS+wChiWl4hT0wsQOBGExKztymbdIlpLGVHp7PzZ
1kALgylpKi6ylpIQBxoDWZ9OFsolkVRImc53octO7xWkL3v3hs2s7TbsOFAbdeEY
Sv0sFAzM4z2FaMZCR/xFD6bZ4fR14UwdPSIyZ8TqIPFeVbYah2kLD0vi57GhAQr6
n+OsU0ZHPh4niJ7f/swbm/G6q4zct2gFCal3Qn5toGv1s0oRe5WFmGn0zltDwCDm
6CudB0PEONMnNMazlVuIkc2ikWptk4jQP0Y87q6Iy6X1H7yOakmlx3j0Y3VsyTLu
cOxUYFA2itHXu8w6uMHUIg5WvZI4SQmHEw3ASZjrb7tTrE9A5MRPzr0iF92TajbO
mYibTIfzeLPAzN+tOP7KUkNKa0KwmpePuoOFYOKGB+tZeWPbBcFhtntMexF0Zi8p
2YKcJBSTwR4QL30CkZqexeHJWYW2E+tyDNh46mRVN275YJlbK69deWtWvzZe4ADy
rvqyuCCpMiP2l8RB0MlfjLA33InpgSdcicnQCtFcZbN0VKWReHdNhkyjcDHorVhw
MBPk0Thaa5BHO1EaNhn5Dzg2gntcrLOf4kGBO7rQSXrl76V4NiiIAQEWVSuz7+Qq
NA0LQjWMyLfe5MReCmq0lHJLWy7TcLtsytGykjmjLUVURO+edPfK9XJ0GYCnMpZ9
mIUwdFOCZAYKXJcSllLNX+fKIn8JaverpyDKhjt6oEATdONFxEtdGqdYgFphen0F
GpRSE/cC/bZkgwBgNuvdlhoMHBLhSvRLT0Vqd6zZwLQvwbuiKaIIxKSNSah0V33y
xM4wrrItOjubtSLrPBT3Ez8fKrBa0gj36VvK7eGPx6fquYL7G/7wFF/naNyGh929
S6UWTCUAgOslIPYh/1yuU9E4krf23AwckhHTeoBwZ+c8JfsTiaXWr1dYTHSKXkPw
unAK9jw/u2HtlfzGo73vs88WxCXDnMYJMmaidIL6N04dIcWlB0qUab0Dtlmn/qoo
MLxMSJU3aiGArhKSeMXs+FG1xf+4b681FDlxjXl5GqSkxFHzu0rGW9CFTpE8N6VL
AMCk/jsuMTtIHF6uXvCndUckO59ERv/3wKXWVYzRV8V8reUvBYE5+fCAzCT/kZKe
kp7APbihXitc0LVND61ivh+cbU3JABHpJO57UB4vobJffme6MYglcKmbBGgVR5gd
OWxjJuJQUyvhTlwuIS139Vb1x4/YpplFOHI4s03Kk0+aFh0NWXKyR1BSxTtE10Dz
GI8J1q+XGX7n9pIsu+hBYrOglm0FdYbXByvdR7czcgkrtSNvsxLW7oS1mkP27xW7
rpu91lfAbZxbjbyFOEV6bNkzM3PmcJctkE/LfL9oJ0BAE3OzqjIT0p9S6covWQRC
WxPnyWBwEEE1zGVs9VzvpQSiHhA1mxrrbtP9zjzBJnmXdThcoAUMdKTA1+zFzUHp
Qz2qHPNa8gR8i01N1TpvBULxtg3faIQ7qzgYpvYivIc2BhvkhrBpgS1UgWOT/7vu
4vnuyAzceNkhdFL3C8jncKSF6d7CUdAMdAKu0r6GIz7inapXkM0HCw1seYKL/yxe
K01eYOtJSsMrpQzaoxVoc6gQHjs4wZQD1xYYFoLccDBN0ZY/ruzALd9LgwQMN4gG
8pSQUw52mtsIByQmDRLEny1k6xl+liQiA9G+py40k2sEk0J6fwBG1xzbjogXuscT
eBlbVzou+xOmqKagYd3yk2bBreSP2AU4Zdv/mwZz2r2CUifeWIui3FTnXJN18Mm8
x3BiLjC6w1eZe105vMF6R/WETv5cYLSOt9/24XxS4HK07cqPs6IKM7wEhxt9U2BN
iTgjrYaXunMv8eDs1Mdtw4ngROUrDFMYEXF4FCu/GEXd17WmeRdh/+rsXLj4iBcm
sxpA/oj+v3q+g8tRCmlN9lsPzS4aU1EegZePdS/VCIelaC0kmZ6bzd3q8BCxKTQh
Y+4eEvDZoqpH9Mmu8yYSD2ihPC4mfDQlsD2NoJOhc5nCWlO/1XDhI4qkr8NND4cp
+Xxxdfkvg9vfYA/3epnFDbM/J3wWyoa60jsQ9tYjXOIOxj5nf7tvWW9dw3Yn+E4Q
Fi9VD+NdRTuBwi0+VElJcMtO7Q1i/3FUVuSY0ciWY6t+J/QRqyF4LerBaxJ3DaOi
Phz9JPJIX1bZL3jgyhUXCEKSMe0Q8g3Hf5q7FkcpwzV2R1HjXBvgqPwm2517fboL
U/Kd5V658hYweDZi17nyC3pdkb5l04e6EzK7z7g4bJ6wNmlOp2E40tE/LUl/CmW6
IYHwa6bQKMeKWgqEH1C6o1goyJdFC+sqNp1+Z19BDKZlZ8rA4JszlKtKTH2URfHe
5zq0yYNMKAE/FlMYoa5WGq0MkMGzxTGc6V/aURdwEYtEGZ+DPTkyDEfXPvC0dTGG
eYYI3UcVmwxYr3ssRm2nhSInVlwBlZVaf8vojBKP/UtJKXb4DYszEAn69s6MDuym
oJlgGC/JfnABKuPtIR9SmGB3SY73C9YCUeae1ZlZ98PJ45mns/ilA6CbJzUPVS7J
mAKECnxo7aDUqXNYFxHn7dPgvlxBTdQgmWIMPzEidzJH5+gaFafOcbt3UVyH0/Rp
TUfGgsSFCTjJwCQaDNupbWd0XNOMQj9RjzZjjPxgHeRP4ScMMAMRlznzmCyQWuw/
yCwJgMkze6jXu+RxUBazoJL/qmNdnjkqBhqdsNr2VJqWQupyZ6scuEW472N1IY8B
kRQN0+vy50XH3is8YwipDx9QQgjkGAcAkZQh8NzOo0gK68Mgf2c0LWu4WD6xlkvD
LXlqJ1J0qYHMmkQYw8BJ0p79lcJsvDS70Klp05NU8SYg4xhtZwpIgstlqnLIDCQn
lDoYIjBqGfxvGtmh0NnJ+OOoPndpsaR19Bm81yAPP04zXjL/MPysO6SsRAp+aDzC
u+Y5rlxijxxMC3NmIOU6PMKgpv8wOAYWbMdCWEIruuPLf01XEm4l9IBmrdDCEWI8
xAXeycaMMcG5oOlCfFXvTBuMmBCUACOp2DQEr3+lpEMDLvzwc4oQUGHfsQVCADFf
iCKlhVBzWBlQ/QVsFTbieBwT+FzxOHs+DUFvWrSC4I2phN1Ll8Gh0hC4+2tK0E83
QcFfzvrIDOq3cPOBdY41gXd965sdgUkisMEdEfa7DxyYNQFFQoM1WsOuIl1xjm2V
atmj/wbCb7SUGlWUvb39oCEKDwYnCPTqOoxyBiuUeqzTgPaig8uVFHQWvYS6Er5P
Cutym7NSAdQGuw8GjC1Z2I+QPgdHR5BGVqtXPS4ySGFwymHy3dGM1wIXmZ2cLI9i
yCMgMspLc0VpjlmZOoucdLMOodioYUwRPZHCdG6xoDiiu3cnBJG8RyycnDtUOdMW
+TXv35g35tocbyr+KAFvxAAKOkcU5v6MQaFEK9W7WeXe13mS9Ql4H/6NXVjFhxS1
vmtNOoIZJixSDF0euNOUvUFJKArdgpUgzC/BmeQ1iss/ls2A3fgnHinLIGbAsRAF
+CLzUBXJV7h5bAr0on8hT9pRblHGZMnDc/djPm9knO2KkU9XRs1gOVNkT6MAHCTb
DCtwIAPrDlj94WmqQzUHKqiF6KdzPgbWJakMNq8RXXrL1C1R6uicqXqq7Tj+v4p3
iU93vd1GeE8YOR2gyzlPtnJmP+2wTwtAh+4NmrYRsyQ+wHrkIFSsI/tG24Qlqj3E
zjDyXB2Gt+ykdof/AdNisrwIn82ZPalmLTBg+DJRd927B6AFedEw8ExnziB+St9T
6+2Ko9zljLgS9wvOkwG6Dq8iohE4sCPI/u+95vmm25/wy5FwCwi0CK+nHw2+I+Al
CFWraLkGS67z3lATtUjhywcOjuleEG2a/eV0bG/bN+Y+kXIkCUlgJXygu6VAxC6m
Fc+2ia+pjTGCLW+KoMpflPorPO17rQ3nZ4QY9ns04LAvZYWW5PVg25u/cKyN66YC
ieDFTBYt0+ArwQKtOMqPVW4gsSxStsha1GjMSzoWVuaomAYdgJz5aH5myTpyd5Pn
bC6kA3Bd2CFWwTW8vhEPlDsqE9bMKsMngDXQ9pG0MeepX+IRQGsEAIN6LbVAQl0d
EEWLvuAg83k3girBZmrXWIXm5LWvexGt7xUi2on+FeE2HT9AYQyznTBp1YR4LN7s
FHB/pq8A3EfncW5E6oP5WjCWPfeujgM4fvjwR6yMn73vxtBncNeW0N1Dl3VL+z3d
Gm/lX3ViwJBuGNtsx1R4RPuPHGisrtRs7b3viIUqNDaksggx1JQlX2KR9T+P+IJ4
n3QozMUGpj2I4X8qxzw+kwPOpgz1gg337QKpK6+9F+IBDP09WHkCW/nSIBoXLhkJ
LvlBIeCoxXMxE4Ej7X0WrUSnX0re7gZtJMPZctRdtF5oIvbbbhgDantSHnbtkEfR
fpT1WxYgUhjrMUGtQNzPyE/oBFZ9ztKMM6a9viyotAiIEROkmYw47F5iz2n6ovT8
RHciTrgZSpOfMSe/xfuuiNRv6ipuJEHxD5plX9pgxZeZ49FQP1fvG44w8dclTB3T
23SztFoRBObwkUNrIuhPFAEVxvlpjP+hNCNTq7tWh2EvVRGzZ93VjUuVg1lUp7ey
o/4UIagSvlw2TB1lWGNONm6c2xMmoA+FGZ2wfaqOtiDzhtNeBgS4e8GKWffs8KjQ
BtjWmCxE4davYHC1fZz6nQ0J1FHiVoC7Oxey9Zae+Vd/U8rKAcbKwMEWbIv9Df+L
4aLAWJr2zsGNjee9uv46klKwKblv11g6nF7KmiDNm+rAhthmCYxaIDD2Unr4wnvf
qYmUcmHZtDifZIBtF07J8AFH/uZocHxMwx+3TaVDNjoF0mvlMXzkNPEbv8vH3EKe
BKa7lkhmv9ev7DuaMGeeP33Z7c/6vtGJWdfno706IDRjxw6iM0NV435bN04nqX3r
HGht9TkUfaw76FI/iQ1+5gHkm2vrdU6LlG8DAGHdL1MmeT8BDtbnChExHlhrDyd1
RlQtx5UZGCbcF8VqDcHd7MnLBcbnsSs+zLVhAoHXsfagaSkSbNbHBkk+ATc6iIcU
5Hqw0VTsEWFB+MRSFiF886jAc6IHbATuueSIjslnedSGEqCFAqWO4QK9x1OKe2ty
WjIuANqUGCLUnhkSvnEu3aT9EQc8tXqtceDggzSRdXh2c6TfT7AqdWyT6zsl6luz
Jo04/6b8AjK9aV1bcV+HRK7fC+ZNQlLHtbQ+AuW82ZGYkmQ4TQdvLkg1VQubiImJ
CtZm+wNHuUAC0sHJrPFKBc7Aib/zEmcwHxbU3iHi07svU8DA+sTU7uIXTRdB1x9E
MYCJwkKo2OVeSiGTcU33ij71WEwP/MzTbTphfrNrnTmynPmSJiGOx+z2tqyVUta5
I/Zg+VuHPUmQ0QRnAqy9XH1U3YEVq8tYzP8VkiXrOSnPHPARbQ4p8S+ubhp6xFrd
AGfmL4rBndcVfuFMhHtJ/hdP0E7D9A4H5itqkpT5m08qkM6CqjCQV1MFXahHOVZW
GagIPpIfAiiREVGuaygkbAIxvemteLdMve89n25g/rZtWrmaI8RSX69ly1jmJENb
V5GNIQ029LsX2oGN8xhbCrMSfseDjrenNUnUt+54xAYRgZiG02SHyaRPjYiasWBq
BCUJs4bKwVYfyTXZhVKbaJJFyFfWICfdB1CQQhAu12HicF60Y4HRz+N4ftVOHRxK
gq8QcnBHKwb67ZVCnxb4ZQSIzWgSu9C3n3t33RnoquSroFx27OzRFSg6Y2Nn7J9u
x/C7u/abHenmI9roGzvcBBxnhh3k3/v1zigAQWkfBo1QtevBPy0UtLlAJZWRrG1u
++pHy1PqqX0ZFZna7qHsd7fVTdqwx9RIbjEjkaD7v876nO0r0TC/C5enmo8iCIRt
eFsdbt6tICGNJjvT5D1FfcFJbjuyq/MMEREfLjgkzCSQbSEvcbgzGPVgoHLQn4DX
6euZS6plz3jKDR+d45yhSq68UZrHqQyKlWpG5Y+wNViOZlyu/IN1pMw4qdIj7TcV
u6GBO78zYiMSmBPhpd56yYkS3oyNcUa46MfKuHEif+8/8XidFYRF06KblRcgnhm7
B2e4vZFyqLn1Qlc6OMiKlx79qGvUzO5R8clPQzLCR8otRdugCT8k2zlEgQM5eJuU
wcw6xnJMnQ1k8rMi0P5JgXDnCeiy2XMe/LHqmy9BLWjz876h/vGi7b4fvEaZlJII
KWLKwDBGu4o5JdM7qqaGB9U731P7Kqn5uyDi7GSRMRnWzxZBwRbBOk6KlCv4EPH8
wuiBq9xe+ujwrE1LO+OF5EYLHFDDOUv9+gZGUcfz9Uu09iATmFOjJm58D1aNdmQj
Q7kbDI05CU+qMOsaGGuAKnRPAlKAtccSzo2PDlPiChdQ+FcC+q8mXpHJLe21Vpev
udt9B6rQgDm5Yqq3fKmhh9GTCxAc6Hc1py7QSLfc8Jeo2EoStvkrLV5QvEA1MIbu
7WYt+pwwO/L6oorKrb4v3C7ZeoSSoG/WjkN5HWAeHsegQLM55JhxcuGANzOQDdQS
ug6N5VYNaLNaJrRtngR4hoPqYVUhiUeVhTqFGg9yc0t34L94l8BfuVzxUij0g/0I
VCJbryGw5lXyq7vMI1GwoOcHLaRiDBq4+mBXnfJq2Oo4QgRXLksYZ/Emif4pMJ1h
manLKtARtHa4VMbiokIyfLLT6/dw/SRrU7cSucL9/NOjaXc96BS05cxi9NV9hFAW
aXimt8WoMNJRURg6Z7vor//fjxz9NSImDRkYz/3q4FV4U2+RshLc8QsgPQrETmT1
xLIsRKAoN6nBa6XocoHgz6G8XXBFP8wv7qD3HlYFXnrfqwk4wFvDWChvNI1ey+B0
A3aXcbOlbLJwEBp+I5jv6IhiZpzWwMFDopuj0oO5iv527+ymVzxGAfDnVyJe28Dd
DnaK0OkaSrb9QALT4BzQ3LSMLBFBgPbkfsEt9/hkFZ+Dhzd3oZu3/G55BsRaPCrY
o7GOCVZzNUbaW8Tz2j/vRDR8aL1Myw+fWce1jdklLtYrtYX/haxDaSYcrcOuAzqS
M1Ra8trwmAMRlKbZu+Nsj+IB0Av3MhQZcteLOIIYG0DzsPVuYChW02vH23W9wBNr
TKaQSQySTprQ7VGDS+xaKlArNJCB8E2uTB3phP9xVJDE3DaEfvcHWKqSUtYSek7o
OxslrH9fIaysYF5PR42ALTM+zPKVT+yq/2nfSZKjhwA+QnXvQHFjEk1HqWaHkkYc
/sR7xA96junWcCBmPmXlKudThHuB15o9skUiGzvWhBrEBzuvIhDOYP9Fa4/IG3wM
R4ClfUIm9cqPUq+YewrMEOP7LjW1vpasUw5dFAB1b/bO/Zsqk+ZxBoFYWiC3P6cw
ILyQgJBH5rKf36ipugCzYORQWwfm9itK36y9x9q6PpaOToSuNfbFC+6cX1w8JNtq
ixevE0BmrUTTF55nCTWcXZr1fMdtLSM7WFCHeknxE09fsMim57lDyOft1tnBl4nB
jSZLAZqXeJmP/7ahtjggGs9O6Y3wQuZ1zYy/S2d31kH/BiWwh714VkyxqHU9iAUA
YCIcFbbPpRXArhy+VMwqJz8ctuFR4BkfR6eze6g2vJMfy1GUsPw4MjC2Jm7qMZQz
OP7hBYeb4dfhqIXhNKQF/qOU5hvg7+gLiuVVPaDwIYlNmOiXwbtU626AyCYExYtO
1tCm0yBBeER4upXceACx1/XdUf8M0Kkt5r4ZWz6ZUS2dAjhLwvz9u/EkyOjrqlUa
x9nD7zE65zGac52WPT8D9+AaQHtHTfl8KAXxz5dha3XdzJktGVcxwBEGn06lA3l4
6A8cnJ1K6PX1m2aEWiINjGpqAFjjVmJCY45LV6ccF83JxRDo86s0ssbSzed7BDO7
Qkf36o6fmUjlkPAFP/gN80MJJKfPp0bZ1NY1B+Ge8i0KlfmnCJ3z/Injh081yRkc
9MI/0WVjl6ZkrEa76Css2uw8XfXCGVdD19vel4+RHvsnlUaDa5VcqeQJSAc40Yxr
KzM/kyMn88i72L/5zi20yohxIWx7JIIczYjHj0D3Gy9bviwUYtVRU/J2s/FSRZOH
VUcR9RBuC/A3v6dei8wYDe6Zek04S13dtoazTF9P1jF/pcmgIhJuiNMFyotADkDy
QYdY/rYMsFM6C0M+g2OO7wLETOEsARvYXvsGHhl21WscCEC104rZKdd6axB+huF3
YwYK71fXWpAgrbiRmGOefJjGqhcAgxy0JZshz3mVNhWBfH69XPqsuNKPYA0blpjx
NvWfzWbXgVUmYWTo2+6AFhy3FSGeP3b0VpKVLsGNCFdlMQuBA9yWSXT+rjoLFRCZ
2JUlXvVUZzzPeN1RtiwqgAWM8Y7bWo9hX4SROWr8zEtUfEtx7Dd9qLC7U3s9vwG3
w66bGGpcvhfVLS0VWJJqYsoFjsPo+UNs6eq4K2AQ73S+81r/MKJ8hgQXyPpngwS8
8tER/XJgqSqatB8Yfze1Ey6VYZ41kSA56vevIf6DJc6uJTtfbSdCZfBWSy9c12id
wc0psm5XNw0fCSNUDkcEwwfUpzAMWq1hVO1xe+A5tivbkVEGLYOerkZ+uzhvdy/4
M0t6qbbaz55XfkuC5zYyECb15aVkNIpkopKf1huB1D4O9LpeJHwGIhHZXGU3OyhA
TdKDNZGU2NJmXOfUofHtP0ocW76/d5H6mrns9G+0SQbLaYLzY7byF2TnzoVVfJI7
sztysOM7CMvVG8RK60/JCG7yNMaiGkWkdqkrdfkIw66hJqcwzwn+TNA4npkHi3Ss
Utezi8/cNrr2bEZlgkECj6AFZ4QQynC/HB5mwb46s0ibP5MM/63LZdyBjMji7OY+
KVl0mou5qxp7kJhypYbFeiZqe7cnMf1aVoSwMTxeK/VJ83OOhFb6hxN4yxBAIKRU
LFWkLql2iDCvxEiaMwljsffO+VVkoLdeXRSXnbhEFonW4DGTzu12Mp+HQHbYi/uV
y6RUqPHptQNk7D2e0fF9uyGkc2VqycejchZLGbgxSI1cYof3nZUxANq+7LXduL4/
iVmG11BTb1teh0RT7XAbyM4ZGBR9SOvIb1LVR2djS1IXAUKyrRAH5ALQKPPxZhd9
L2t7TJTwI3wttRvu/mV06D8I+wG2VTxZ+F1ROKmWKCi+dtc4H76NjBUo+C3qgWNH
oC9crLtA8nFyxTFwST2GTVU6qWCqiHQF33hDqKN0DzPzX9VvN8cLCcFtSBeKIzB9
CGu2IjUuM0KE2rsyPjYrHtvfmrUxppTAE8xpJAxeNxg811guEimImQ66uaseYzbb
CPA6liEHbSNLrEKIF3llD3g5UnRIgpqlcligWlx9q/X8a4rIIOdOITyZC++2TD3Q
61Bdngdvy2RXGtZm2ihkS8OSAicFTFpHf0XNbVzC3XkvmJNT85qY8SXwYj4ZT1QA
Hu3Z82OQFKk4gwpmfuzHGJnVkX4Uka9xnvZe9tBQNvPy3FjzP6lVcXo0W0CUgW3i
CLS1oa5fAKFR8x/NZy3ad7o4pHxlpTTLjBl1+mrk3G4tFYBBmiFa8W2N1dJ79zCi
RIvdziwSq3Lc4HUkpjAI1HGlI/p2ld1DlmkzyjOfUFdfxVWQrTPeIQUlVhDVrkac
PwJgHPub5/xbjdQRWTEQL24L/loPeq7+ZQl+ouZFbb2ZIAv3AQQbsOkGroANEWlI
MR1MX2SKo+144/iCc09gOTL1w6a5oalSBLN+bk2pizaxmcbg0YBS83wGV4kAEXKa
gVCLJb6BKJZB/iJfC6NzbjWNqj4s0SA0DEdMfof1x/8SKW160N8u+0EQ4Dnc8yDb
7nW1pxoNUsGT5vAM7niaZXTm9DtIRCAr7l8tJitG4ov+ambm3JgLEnenh1FAxMFg
nOd9j6P3oWGX9MYzs1MonCwxpKzTe0lYYVH6AczDjItfIT6mgL667WbcLd5k+KZ8
arHrQq/+CMOu5R11hH3nZk5WwjWCtng4yN6ZBICITi1Va2VcsS8tbmyxrT43kaPr
xMtTwQzhYIUvuIM7kwfNmjTZIm38gCHJUNpEpig4XaY6Y3vPSbQ0iKHblIFDUfmB
BgE3b+Lleq1dqCBAg+MtThLWGed1C8Ge9HZucTfzn0SJKEaE1mKBLP4g9x3/ItE6
m1q8QmJtCSuEZN7RMg/lgp4dY0TvpcKTY5ZKTWDKyyyRhGnczPPwvVZX9n2X/1hj
bPohbAKHPnZhVnunFuDKi58avrgATDssdhZGBs/I7Nkc0PR0DiJhMCQ5T/OZLGoz
00dncjCnEoL9ILxGSki4RN9PACpN8gNe9ARjXjACUy7dw6xMda5rtk6aDQtgQJVp
iB7P12uanbNPiQBlg89GM/Oyo1RwppfrXSCy3hiEN6KmvKj/XbVF8z0o110kQ/CV
vo3M/1fJaDOZCvWBMyOs2Tjm5J902SxgkVb8HoZIFBbobrMc7QlxfwXbr/+8eLTM
RYuGGE7zF5SKSwF7rWVe3u+z1MySCkNIXIY/WkstuD1/2S1yLMfDq5z0iVf22kvR
V/JYM4FcVR6t/fXDGVa2p3Fdj1SlVxIgbdpT/AnU3zli1CThGdWs1Oab/aINvDD8
RkmYh0smLHPsZqL3WqcX7drrLls7Os+tBw5EjgwliHmWxApAf+eUefTMtT03ds5T
jLYNM+cDB8uehDOt2AanVIsMfM5F+n42loJg713HHFiASf9t79Ua0CwqCoQSDK5O
2clvsbHJ334s4yOG5ItOfYn8BgLWxxAUqmgXYcUFCdT8kQY+2Rgc21txYhWA8bId
vJbQJe5ydCCVkAyzAmgq4PUDPvQP5wFg007Iq3Y95K3ZschWWzmRIFaILZsFMH0D
JmnOVmDVsOKS1ahNVk6Pwwalqa+McS3ZQf5OOp21PGVMYq7C3Ak3aC5q6HET3nmx
MBuaPSgrNqzUdcVivcL7VXXbtrcqDOvoLyAtxAfZrdapv62uz8oy+fv5zARvMLO3
sRbeiQ3fselWSyDsYlD5OO1EwVPLWDgQemSTwVW1yPao92F8Emvo+DqqhZxci+Lr
eAH746FObH1VY3Vf4odBOFV/oAUiapfWrtIzFCsU0tyFFQXAyZoXa3eNmefhen9G
a5hJZ/38KII+vIDISp/Vainss4U1TyLOeypOP44RiqCSG3bHeeVtgFAnThM0p2x3
l0L9z+ReDkJvyJ6E/b2F4lDNlr1kvg+Mmi+nJipQZqRccK4irE2jIq1DOOh5gCmF
gNtZdR2tEn4wD3aUj4poEg26eKhRlvTHTFX91npxarLh/OuzqyD8ABTlIdrqiCWz
/3xwVNYDQC0CD5aN5nsuHAYhA2SpBFYl1ylbOpo+jDzRcyYIpqimAg6rqqNAkNye
A599vUwthTSmBXDicAsg3tKjs4NxFnZzT8DEIkYrVLuOmTRBC5VzTV9ilJmp43Bu
VBX6oOJh99vK3Fry7dh0RwPlaWLTQw6Kf9lL1/ykSsEugykEJexlKY+RbrLAZ9tn
EZBfoqZG0vcTic1PZzmayjPMv//0WcL3JV41Z+W73nicbOSQC4PgLxLEHFbERKN1
P55cHztd/9ps+sjh4eAYiXIEOTymCyLVTAc0bBFkcRVc4oNGotHgPqVszFM8wS39
qTMDHSsbMsr+ws7y9gS9gB0RPynoLQDMzeiZjBcCQUlOKA+loxdxkMlJQ8IWDEOr
niuu1ZpGMdW4ibC++PjyJq7BRAwaxzJ/KPyU8dsgxUMgxS3zK5XaSNvTRVbB6+aY
srjz6uqvaqtWoU+umbnR/a6HCvx7E2BiY5OYiAgkiXGoT8xIt4sfSXl3D0buhVOy
wOm5ulH5C78bwZZmN4Z8MUyChrWZyofPv4IjK5JfJ4r8yFKGTFUdh8rIAX8kkzfW
Eifb5GqbzI6Y69H513fSjJ8ndxNJeNhT5q/f0cU2EDOynFNmVfnXVINxq8T28jRZ
88RXK0aQ2UVPr14M/IXv5FNn+vDr4A9tZkjmQygzlVeXNPRhxkB1Ws8HHBbidnn2
skQvGEhPeSFIiJtu+w/m09Hc9qAuO6mmF9UbeLBXDy/cpfLEgHwgWqzPt8PGd5pc
fpzOVYd4iYpNdD7vZglyGFC3vXAEidkl3TdiaFGTsDe16fZnKvsZsnfFGpZcDn0P
CFwGONQw3WYRuAbgFaXuzpmEt86zM0PnHn9Lv+JdsnYerOF9LzlQ2Ic4avoJvWhP
DVtNaqpOJ8ClIpldWjcwNVux4ZqwUcEfHTKW5L8LksQnkGKk7fRE/65sbYSRKaSZ
6zXHNERbm2S66UuQQ9dGMl3eVWKypOB2GO5mdBywH/RCyk5c1uXs7BuJi+eS+A8K
dkinMqrynTEbEX25jTDCRFGDUQ4xeVWWK+sFPbJ060Eb5HsS4tu4yEmcwFtqotT3
BUy2JjnaWSlcY7yTo5OFEwdwtKq5Wg4rAB1R5H2uPY/IM+Hm0YDtBQ53jJ6NKolO
S0FB54EUafHU31FEFC15gcFWBSTGPvxLeKxi+vdTcLxYnKUk64jb/YubzSs9M6ou
6uqh4uauY51pkFHz5XJlhy+8msKczUVvXpAVcPnp/tYP3C2xy4MICDuSV4KCi99k
4ZhqlPoHGVdHs5Fel7iwfXmIg4CZGN39C6LesUSnp37zP0wWNuyTqkbgVKnEXF1K
wZVf9J3um6LD0Rxd+uPYlOa8AMrwk40kEuhXby99HhoBJZkxAt1w+PiAhUDYx+tv
OBB1PQhge8wLk7jnayvAM+gzIS59YRBXNtPDhYR/77v4DTquEis6XQGI99sGsuQF
fxO5Z5E9S9ropc4T9EnDkDhGj6hSUiNwca3ysLlyGUgrGPS7VPSpveP1tSzL2VPm
uFUXr/siPRAS0jMvR3HncDZOx0mYZuZ5rzpR+WACUA3Z4g4Hs9REeJj7k4bUEDQv
eHrB8NGmQ5rxf9L0wrTwN1awCGTAiZVOpeX02Pnj+ogAl4SoZc15rs5DawF70JYp
lWGe/2bmm3kpsPuedstgyoen0WtGb+oCcIObbPvYlxdf40pmYJaW5mjsnu2ICCg+
64ESEp6jML27etgrS75kes4AocvBkaZRaRXrW5Q7MRO18Q28TTqN3CTSnH4DKAiz
AL/QjNAhUDND7D4zzxf6d14vJoiKcn24XTlO4Y0+MIOgbMh1vRYRNfdt1cy1QIz0
5ISB4Qg01J52SqOXTuh0LRpTSeBA+Rj7nqswE2rgngJeCYuSUK9McHcojaOlbHPb
qr4HxwOEarx9bH1mxbCRvY6H/umQWSSumYmpvv8fyx2YZZoDVFLd0vu2gt60JmNo
KbjpgyouvFunTqWlCRvrmmAJsueaJD3JYV8kDxk8UagYBYUmg1ALisNnCX9uH93Q
zza7277ey+9cmMJ0vz+eGw71FQz8g36q+FSoT3IICgd8/fOdj8vQnybF953iCFER
2U43/LLspC7cOTFyFYLtJu3nFQqf8R83cFFgjMdSPC69hmwSLiFZd+PO22H1jn9K
Uh05o3Ltm1ZFSQ4DpwvmSeePZ9IPRssEwdCPvZ8ZO6Zzd0k4erwVuxHS6W2P0C6O
N2O/Lh/RJMuU1wEAy4/2VgHkeQzhtwp0aJoIq+0TfuRaBoybo2IDc88eKQ7jvOEE
hCp0y2SXFyZWctxCJxgjsPrwn9ZO/PrxQpsQ7tpuN77G1M7uBUBjhlH4YghenHSu
7MR3uK3+K5yQ3Gc4niZATU+9/tcB1E7ceBDBs6eMUwdb+gyhaZ149usemxNE9cHK
IFv7c62gL2NqPqxCX04YMC9uMwH1ARtTlJ4P1BLh53TS0HsESOJV6iMVExfu8akm
Vwpz+b7U8Cge/EUgrf4UgObIFXkmFLS+wjF1EySaPvsevgj2qr4Hv5U/jYDO0MfE
PHs3+YKUYeu5twr91RgpESedHV+JF66gPaKZGFrblujbfaaqKvcLWg6ALKViiw02
tkSPMWNOPHLCF+3X8w+5vxHeUfrlUb+i7onohG4GRtX84rx9Cb4/awncoE8OCFSQ
FJnQmtuj+3//j8O/uUTLNjNMwYzcdhVdDt5//z4MmHTsfgrWv3gBeECZhl16NqED
q0jY5TM2MR81jx4neGlT7x222qtqS7b5IlY/JCa5Q081HRL/hIYjCNzpuDVZT/7g
8ioJ+05G5SfI2BDjfnRUBdyoOCtY2QuLUkwtW35G1QcwN2n4MqfS6baYoEhKaAz+
bVxGWCBg9jzGF7K8akypWWbJnQfTkAhzzemZgoxeoZBeaztXz3rQWYXN337WHdX+
KHPrdNIyJB39mCt5M6XyRZwE66bR5kmHVJD3GHNSMH2w3huCHKc1LQ8GAvBt8Cgp
2edve0/M3l+WjU0QurCC5+H3b57UTjsVdghf4ZhFzlBi6Iup6foCVtV2rDqVzNvp
2A8ZL6ZEL3XxQXyy+HN9tA/IXrrX9iH7kEUa+krJQi7H9e+/8WvBzDNW5zgd0od1
WPlgc+vvtgnB5jqsRg6kdAwV/X6tq7aSmlJRaInB8qXNsjYtXDtRT4h+T7olxrEI
gSnWmzt9FYsdDczSXF+BxOUQeIg/b1PGGkq6DpZ3y2djs965mNhZcH9kZ863fDTB
SqNdOU6H3w3IG63QQ+l8EgzfWKHfhlC9p293bx/2wAKzemfTLBf7HsQo+88tGtdK
36uV6sgWZtlVTk7ItYsYpbT2Iu/FzRv558vs/HdQNpEmx+4C/fBE198tnVDIgyde
Y8P5oQt8oMZzj1MkGbWCqcKTWeuiy1DRA5mrSmneEwbQeAEPN6pI4XHSXT9dIQt0
9m+lrhBowmgI/LunDHujri0jAtd853oSjDDm6HYrLjCSaIgK0HbWKcSub6bFbJjY
r5JVCSwyjP5Z9fQI2LlRdER8egIgsZLAqFnKuniRCDrgUZ+ukzH+qCQRsnAJeeOy
6EAFIaMkmf3nDNaY/7wVlntD125mTvXid01yI3/gN9WBcGTzRZv7fzmVdpB0NenR
9Nhh9dc2XvJGexAL4YIYUvFK7hNesGu/9KDydoMB/enUBigh91VQ9Ss1NrsUoxgJ
qtvnhz0DvFV8MMHdf/T3fEq3mbp7wOeR2g1LiXFSQpbVPu1xKQeCfl/QgREtZ6wt
0uRjPj0Wssui4pC/ooeHMOW/JcnR1HZFEnrS0hu5EBy1OTyPMyQLmx7MIXisLQeZ
fggNElDe/A2rwt5RzeuSTSWsA1/2q/lhfjKBI/dBZipNUDaualVRqbNWJRH10wjx
jBMFe57ei+CvLmER3hXOEoftNrzes4ZltnnRn5OCCmyk8Piey+PtkRhNJGA70WFx
x/CkZKz4WeXqOJtllKoFVoPuwempaoppoN+P9+U0jvBQzq/mIvvjXaMKdinQ5lG4
9wuV76mlLVCzCJBlanOdLmO9yocyCn+kW9prSTAaPD5T1dB41wTjp7GA5zCo3fOZ
hpkoLlkr+aSRAWR+hr9cB/534j+7qXwyTnqF1Djv/JwfdrXI8fCDR2thlrQcSAig
ZcLyyFIkM0ONV3ILJJyAntHnr9Ogm/kq/PVmxq/Hn8YFtQrqqgpYHZYeP8SqiBkQ
CSIPxp2TFcwqA+z1wrd550rHSiNWkje60gc0bzLcI3OiBX/BOuMp/jKE5F/ucp1U
oORsc8QNUWNQKGektZ8nF6wqbi0W5NaB9eYiqKSp49B/MLTfq1vsvRsLIJVKl5kF
2ji8sXOlyvp40fd6jMsLMhbuSuWqZLm5FSGt9bk7yBm6S9Pu5TRCI0tIEHJdUQUy
yWYcoTirTiiHLeEroOTNiuFLegAuGKKZya6lYO7TCR1DGajKx6mES13Zsox6gv4q
6gqHAtRPT9oGVenxxuHFMdDjer59kROXa8pJ4nJQdA8YPqNU0eM8MDUZ7UeM7rFL
wYDZVVd/Dvuku38MUOCTzjOJrp9wAU/7rYDZqo63JX3rF14Sv6HLdXx/HAj/gJFr
Pxf3vGuLd0Hlze1hnpdz1G8p3wgEsMnfOS6ZmETMHQedAv9Y+KOOVksfzehHywxA
MuXyvCpocTUNdU5dGqIuGG+Zf4fEtt4V6ekGA+fsg+99bPz3NPqQenQkknsv/gAs
AqnQjC6leNxr/1fjGMcjs4owQxeNg+dgQVsBIVY2xr6t7NqkM7FPBvfO3C13hFax
C5LTkeBCzCcJlsmD5AHH9Vimi51WJkpmTxS/5uWwfttX3O1D471+enQ0xQdQwces
AVMtoK2/IGSlXbbanE3h3U0xS0BBYV/6QqaWUNz6eEbON6Ofiw8mwZhujo+/Motz
wxwHGqT2zgrzwI2ZALjX1vx5wuXZSVrMyhprc0nU7qO58va9A/KWlAVXzofM5V9/
bDCrZIb+3APk1qyf1zIrcuuDi4WzpFBJh8+a7f7QfmfVpnU+6TpvgqmXl89ql2tz
Vt8P0eQ1r+sKIenYBoQnS+xU3z+Y02GZdLcyCKHY8hxqurGta0hxP7H8kRSNgp3k
VxJ5yXwOXXz6SvXm57vSsf97VTRPhRA7YuzOOOyrdX0HMyx2F7dgmbiMz5mYnf1d
WoCMQ0LHRVnp36IhuFIVeKsoJX9yMjDMHzhqfm8ArYoHwV3fMFv20RVcmgFW1D+k
eNdQx4JSEZAIfVIZXNlbPTh9Ymyp3OhIFrwspXRQ0pPXuwiBLo8PFYGKI0Sbahu/
JVdGQBi3sh0vsToNaUnYkYMo0z4vNVRIheo0/VbdhsNn/R41zKQq9RDD5q3UJLEe
yxK4WUomxI3vBiw6Zh5uLb2/FmBGrtMNnALLh7FgD2zcJPBwutuHl/fW7VA7eY3s
inRyU1EO/77GA9Ycd9+GpOs/Xqe6lqxBAeAj+AFZ37FIkcws4AgMbpRSUiMAskDH
8JvLDoyA7+hdqXKeYTUszadlNfbw8Ah5GBN8l3jli1vHgEUpcx0DouzPOFgNTPro
PIuDsLucV/3W7d/JREVsgKCNhDO8F26muwU9qZDGHt17ORb2NSd/vlTYHddKf9Qi
JPYp+jPcWPfc7oTOVCBqBkX1Ngpqhvrk6ge7InGU57kTzaeuPiuh0B+MLfq8LUre
ChWat4eS6bGHHvBaFwNCR5dCPrYkxT9zHC4a3Q4XZK9y0edoRgTyWslv0MLiGfR4
gHlJOcMyWpC4KLlhMzDMS7C05YwCr3Waj/PRh9yPULwHVq9krkPCvDkrQb4JWx+S
oUGWMc6PlIjoo/6wSK/kBVlIA0OO/jlc9K5XmjDWOSNanjfcOfQlJgb4x42z+nw2
EoeMQEzeCX8WqYsArdgW/3XLY6Zs5ORhIq9Q/avxN9H4V1cDUPpLbhNzLaiMSr0+
IuMej0vdbMHHSVxSpGQAfcH42n/O4EV/4+PO41Lbf484u0Q/Qz5qc+ftcR9rx3Wk
K3wMXA89QNH/2FKCgvjb0MWHagdZl11aWp08XM5YKj6L5Ha6NY9X4VnFJGV5JHqw
vTM2XC/kZLZCPecxM2H8O9d5+xBdugmO5NIDnY/IgZ1nnGUeOTas6pvh+VrFx9dO
yf+4d1ZES7oS2Naw6bzrRv/XZE4nYY3EEoMiOGsyYq9kWVz3y50sTeIBF+s9KvRK
ODksKcgNNH8f5E6twVx+avTmN46LOubjtXHbWqOuftFtsC3nr4eaoiZxIDwFqSt1
1rQjyHXuqvNsb/mJoGzPQKRnNkImFo0FjZ9lgDST9i46sztJmdv55+hNd01oFOVr
LkMMCjPSzY8Pfh0W65lKWv1nRcQOIe59uNWXCy3zyIwvu5tIuMHmZXb7nSv3RhdN
fqxJGyQp64jEu9xTAD+jKjg2oCcpxXSXwaeQajwTiTFGTIZPyc885OgOkCvsZCsu
UUmb83oneQh4eunw6PIEPUrW6mjb/m/EC+VQvB+9TzZGjd711hiP9u/d508iG0kc
ILBUxi9yczfQvxzdCIsiR1/cO4L13doAw5jS0Iw4QEI8sjp55pHVCHD9x9eexl0w
CnDDV9jEO/o0toCth0mHDbuu6Cw7U4Cavs5SR9fehdOmYxMI4s2iZteIPwpyYwSX
pct0mQ65Dqg8pgnO7NnRKAM6GDIFCkXmi2XrxNAiQ4yXi1vx5LYQmOcTuh4gQuEd
3CkzNLvTHLE0s/ShBg2nzUDyELll0rGFIJp+h9DRB0TIPzMJGQYC/mW7N3qkJgNR
Pwnmzpz81dqwQZMrWCwmip/mvQ0D7XJdSovtnFtWKfpvdXztfL//raOwRFsu+n0d
asSMiE58Z4aCembv8AKWjQVtullbZH6DgnT0QpAnER6TcjLgsW40DMc5SPFdGHZZ
UgtJ9xROUcc56iP91ClotOX54bktuuL7CJcPz01yTdRIgK8oJbrh8vfnYFnNceUH
Fij4W4SxtfeD9pyakgyMAi0ut2RSx97RlXB83jc3z+85ji6omfJ4wDfMH02T4hYZ
l3NaPyo2gjnxeHxQAW3BbpagxDmxHzd48XKBeur4V78f2u/vEagTwxCR/N7DjElz
YcuyTH1Mb8m50NodTs5Y/9ycl9hFmKUBn+lsDcOStyNRw+9K4I9oe90BLaE1PbsV
9+tvlfG6J9DojgDHghBop8YebWR7JG8iOW6zGboR84IrO6aGk/cKlHsUULh692lZ
vKAAMV1ll9pkgzLeCsipDoWjEBaSdarRMos03a8Qmw29Nl+11dRXVEjyR+16dJRO
6+Q7cW7YWqovDicazk1BpqNhSOAT4LB8VYIO/sxiFtWGd83bZ0aXbAKU7WKvaJa6
WiqxNTUxqUTe7IUPR+pYJY9NaUCN8JmmhY4IXuf5Qjw5O54UmKPYXM3vGGu98peP
v5fB3IEz6ZQm24fFFCHEL531PiQu07oQr68z1241H1xeD18Ne7UKN6H56rXmOOh0
smBH2jDwZnoEZUUxOoVEDVU2TErS3cB2SAtVMEFxC4YplNc8OjIhKJfNk33xzhlP
fPKu9tqlnYKm6UQahZ9NBI7TvxU+bPCaUz0chFa4tjdI9DEryPgh6ZgohbcC8wzQ
7u/zbxEODEk8SHSVmdx3Kmt8XGJ1imKyHZRRV8/wybvaLgD6zglKH0TDrAMs3pvn
h67DngYJE/u3CwWXepyvTJaj5QBU3+5VFFqDxPSdXmKKa6Qjtw122kZ+bzHJHdwu
t0atBfjeDB9kZ4qk4+sURLZVQKQcZ2SQCaoHBpmwUMML1jCPLIXb6MKUkmERFvw7
KNUIZyThKGZnxyApyA10onqRqJZuOu+WBlpHDVzsl4T74ymkPd3Qw226D0mv9rrN
LIT8MHwM0ecojxKdOCo++gNzNtzujIJXX221m1ilkrY13XTnwSmvSypUz0EBMuRj
ec9YvODhBBXMu4TLrBZccbpcJcp93EXVfs4VlaOdWoIYHrp+TNtsIv6Gj2jylvYq
Y4fMNnJhOSq15VPx1wVMHzceGZXtOvst1EzHNRisY46w1WkUcQNGifiQiJ3wk+PG
CSMmFpjevBbvdOZ642m+239L/WArZKiJ551JlgB2ooX05g1LWW7tKUw9b64NzoK0
tldNZOp9W9dYbYLQ+rhXGg0OFlIBnFIib5coCkWvP2iT8vXi6vPqYJi/BVPRifGP
p9Ed0fkocXjjezq2u2V20IUt963yE5jV8mkNCDyH1WIR+K4Uy5Z2Izk7XIP04Ez7
hAkbXvyKIUEdNFwe/ohff9I07g3NMDcSsosFrLnAYChLhExCeo9KCQJdjIF0Xr8E
mxOF24oKYqmXH50KaWJ7W4dVyF1nZxzp2f04yO8l4aOTLM36HI73YXjhPd5LJpqd
JrPob7YjXOihkMhYgtsbgKTFKo5kFtiSWs7kMLRpGRZO5+LutEXgUqPk80KQOpNe
zNWSJu9zUd8uVxiGhZIxRPSCkfS/SbPxy/97ifWTiuMoANtuQKwy2VRM8YtG9f6p
FsBI+ll3g3jiPTxpBu1RvF4KH9cV+FMR9ZDcEe/hTz7NA8xx5mx40jUUHPyZSlre
5gBPz6AunloWu53h3lCSXhv91ELXI2q9y/fMwAcR5QoBuJS7/JxyruCMjoBZq/9p
xl71Zz5AzHgu4b9UyfG/4TFryVGEQBQSQNdhlLh+akW8HJKPugu/+mwrjeAtmv7V
edLL4N/Bgvbba6xwezYM88d1L1Ai7D3nTQ9Q8eOsAmhKTihcbMjbI3Iep0uOuyD9
X3+S8YrbOHHa+j05H+8/ZHQXXRGXzy02zq53+QOmM+PnL+td3RtphYNgc9VpPiZ5
uerDj+UwAJD0GhKlSRr5VuySVdMNfVRHMZZ5Drfx48KUzvQ0vcQ7A7D9Wnys4LaZ
mt970HqTN3SkglMyzBOzCl70rUGQNtjKnTy4/RzcPaaw0C7TK9HZ9uwYmpB7w65E
BpIGi5wJHAGpritSuX+s72qS50UHXmPJHeE+3AGrNROO1j/+ImRokMufa+WjeOhZ
CF1yJZ8b4gOGvLTDeIeBIKSy00rv2RJPQqmJKvHawOO6AKO5SbFLCfpY8iz4w2aZ
7/DRQAACexqPOOjs0xG+Px2f1XQsKs7eu9q9LcpIjukaxbAoNdHzICqs+Oyi+RMV
zV5p3c8QEb4w9EhUkPhgGE01lglaY8BjUHvOjaRN1Vw/EpPWLsX5io3IOEa4ONPQ
I3hP3aEZ0Maqy6LJ/JS1yrkMPXC2WIx4nZHtQWbRT2DDbwOhS7RDzLsZnx/TRLD2
m3It5hBye4/remDnKUr0nSCuGIfXc2h06tWph4DdJL5pMaVpgUvve/yDc0ipRQf8
ShcXiqdhE0mLBuVfmOqH3pfXddyps6CZ8/awcKbGxhVkIjJC4fxE4YuSSbl9C1mz
eKhwJGMyhUBPk71aQYbh7IJ8+EULiSP6dPRh+h3lvF0Nin/TgeWHY3w74pYxzmx2
8I3P9o4/VeqmWMCiH4FKJ4qnfFUD+/iSH1kAyDLz2SHYBNny2r6IK6ExyUsct+2X
wgnlEpcoa7aBmOtwNkkUeCsv3ycRsvJ8Dcgxw+bUfu/q6VhSG/ws1dHPS4wxF4Ih
A6qDgSUA8z72nHosMea19qEdUgJAeEoxb47uaH29O5lJqeqSkeF9MebFGDf1LsE8
W7hLcQLcPfAyKmKbQkXLNrBomT52IZh0vMU7RbS9SBDZ2LvGyxuPpNN0tHjMrnVv
20td369VqRpAbX4GVyzvwQ1AfkqZZgw+ZdmNDO1wHL8SGctFID+EMtNY2bdDWMv1
GMfR803OY70nHkIa4++lvpcfACSl1029eHFOL5VuE0dU2p+Lfc6aDfO7zeE9pBAi
7A5PRnGwkXlR/FnjDxxGafs1vEgLMoh7OQD0bKVbwvklGDh7vQ25gUxN/B3g8h4V
dja7+ueIReIKuecepfsXuSac7IlEFDc6iPaM2Vw5IsDvi4xEhKPXSfYsXCljbIRu
YQuZAM1FgA/V35WMaoZjj3RwKLKWUIFbG0LDPXN+wiwGRKrqJCFBMJGPe/vX80UE
P1mCyP4EyIj0eD/yGt4xRJzLc6tuvl+12TAh/3KkkPW4PxbRR2hFqmmCcJNhu/81
RZ4TpAz9pFx9adRF74Dyv0+Kxi2zmSZwiNTDDLOxuj5x0/PYDd3Adkycw/oeFjGa
goQp4embgAHKYA6MfDPQBADuRurkNTmhZEmVWpC9DAN8N5z7Ei6W6seMt5T+MBKL
0AnCvPpZZnrZtpqQ0IGsSSLgsCP1i8F3w1rSaJoha1T+ozO7b2QRrWqcKZFXo1Dr
xZvraCjnXn2ExXM6glrBaGpEuFpNbBIswzwiaueN/q2i7DdGQZpxd8Vd74uMumzr
yQ6cCWLGdQySiDsldMZFg1OeAlMJlqNh4VTKlLWkqqZ+TjreS3590BWtg4yFy1Hv
VgW7FsufvzX17pTAeAFoeUnmvdFPJIKz/ifWaUmmfbkDZBihIig9dbwaol/Jc5jW
xMIVKMXDyS3ORvs+qFuH20B2QtoZ/zRTLY4X+TvrlkvVqnEfOnhVpYJflXgc44Fz
Z/dmpdpDkFHfXfUhjepJJIljk7eKyNZ535wSZAecsd/NYSSJwejb7wnpFkBLqsK+
8KLN+ytC1ESznJLLq5h61Sa3bhZW/3K2o9/BATGehbe0WB+gnR/3NxE8SHbsvRT2
MsT9n+8M1UNjyr0MK1ZapZASyoCA9RYUy0Uio2njw/Bp3fphzmEhCIJutN3PxFvF
abUUtWabsdWkXB1t+jY6AoU09k6lAVPDduCQd2570ekH0F1EeMx//XgEbJRoESpA
9C1CSybmaw6JMiqbDaeyhIw9PH+6WYzQlyRtC+QoJcWwL/7iVXReKG3kZXWk//De
BdbVsdmBY6yE8AkdW1zBaohfTW8F6DamNCf1FC7RkINgT3rBfpsluwZ3t3xUVPQD
c+/WIW5D17OH0Dh2wP4JH+9oDokQOue7LrAWUyO4rGAEWomoJoPWE832WAospiYc
XG3CdPp8qzqDA6/Rt3QsuzLXOCm/rtHXHT0y9iUpMN4xyiuoPwjZJUk2t5boE8lU
NRte4p3/vOj2XOkPjsgxYLE9rg8CtCEW7CNAIjON6pmqNDtu1YslDFoBanUkSv9j
HgO6DpEoB4+ot7Csf2tMf+JwP094oV0+1dv9oaBJhqCkLvC+1SqzRtS44nhHEtGl
F1/zvyKi20lJ/JHL8PpupmbTzQS8oUOsoViy52jpJDiLEd9sW0nu9NySw9ExsdZF
AfEx/TUmgXBfcwKaSJilnN6AAvTz1V4MM+82YvNVdOPTlUHNb7yCRXw3qLj1EQRW
JysdNj8a28UuTX+W0MCF/NkT5+pKJN5Cockm9ErHGwX6v/ZkLkTk6/7IUqkUv/eK
MZYI/vsdTFpLAtQVEbmwl2QwjM0wbdCGwCvHXTUvlgOZlQ/NJPGv/8JV837fz1y7
LqjR4thYSyLkYwP+fl57GFtyehWrcypgFGoprITRw1C9A0ogWLQ/evwf0AFJfzvx
mK+GzVOE8qkRv2LXf3UQaeQvdrhWPTgBckUEj9p9smO+xLxp7qt+Zpx3BVDqtkOS
bGjPBjivApDZyiunb9Mzmi7zpAkcl3YJg4PoZCP1wU3jaelKK8OFIpsguQA7el1v
FIYPK6vXM8Fdo9Uqak1rDpX5ZQ7Ai6vwxKyELnRQ4hAN9557uO7bcbrTlbT8Qs2q
uH+UaSLrm6GiwdPK755eGRaM26BEmrQqIk07eXmU3TtaMUjK9E6hjXMutFU49/R7
mDqLTWkwPmU1zX061uRIlAz66QHzZAwxB4fp/trZDX7hASUlmrZOls2cV8+VgWuF
euvrHI/QottCZVrsxzmGksiS9aN59nFlZndXAwe4WD/z9ic9jEOugHJpqTOZgK8z
076ul1xMTws+P+awjMGG6vvDmtQ5URuXjQ+2C+6HZYH++T+RMJJDFMxqWv2Tlx70
Lw5qhpC4npjVNO+cRbrJi6MGdHQVL24s9vy+u0i+DIaBXpHxuo1cHTxCCYFrydKj
g18kNZnfl2X92sHeceX3Ca/CnH3jBH4YRuFDJO2I/5+hLbpWS+TqJGdWiIuQYq64
5mTscmZOLwA7XrtO/BTFo9/Odrm+cjZpViT3B70L+jjEcSrK1QQX/GL1Hys/uDtT
FazBXJLFw1Lx9mIqGrMqO2XRcNtjZkX0c47qQS8fh1STYv3PL17riIcLZPIBwVOB
DXK4nWUm1T1CZvRVl1815HDLrBpaKZ5nl+dBK3B3hCdBvKX8KHfOVy0nmNGr9CrQ
i4z44LsOeqFaq3UgtBWuHB6fKluDW3xJ+ji4zLuun6g7h/uMHbTTYM80l0qZBq4n
3F9bCSdr6y9fey2eVW6G58MgELO1ptFAkCYwMAbDZzlYhtdpecNFLwA3SqkX0cNZ
3PyJYSh6+wcfuvWzsv3ns8UetzmBeHChWJcQVE01ZhH3L3jJiP3hkulIw1Xj6vaP
f8Vsy8Y0tXlqTHKg6QQK+sWlLroIStp+ux6jgRV5BMgnG626Zl/wN7qo6jF4yuQo
kHnQ1PMen5khtp/g8wxi5m8OJ1mwSZDxRNp2wCZxBRa1zWdQneMp4/9nzM74OmT9
dRZ83qVTV4933iODEhSEl8rgy8om1kTk9RHEMrvFcRhHeJsnOubVh1mW5GhcWk1n
EZwiKmTyLVjzmsCgDgog2ngKC2wfZAlhyZLZQbvHEWuOfJAzmswiR5YyND+fvPMD
P8vaujv/Ne5eDGmpNGfTkyPj7drr/Ll+crTReDqWXV49HbcUHNPmxVn+RSJKvUf6
C+jOJcF2wzrH0TwxBeoBobsiB/P2h/uSpNXGglQAxr2ipoXxvbm/ABcataDzZiBP
LuxQ/6i7igLUxRqIHBn2kbkIwbEDTEJXhTZkd2hmLbB4xWAHYv0701a32xpwD7v+
1wQuabOxVWL7PF6IiOPT+SEKYgpqTt1bBXGTqBFlG9+PLlFEIriG+ur0Q6rdjv67
SfIDgURYnkDCogfK9QnTj815JwmtOa1sZ3X3SrNpprgAm+W31CsakW/wYgLtGLtl
VzUhYM2+mvVQaWmMGUlgeCwK2xa5DtFrK1yuZmY8/QQdQNYnKaQeJ+Mb3gvdynK+
SO6YIBhwT1UZPIyVZGo2kTfTKr6a2mZD4AAVEyOiO5zcrW/Cuemnvc4YBAgJ+U4g
/Q6DBxzmVKn7s0esBbLC4dU4r18+IX3S5fAsMP9cnFyPUG5kD0KIMys2XdKy6bPO
DfSTOsFWrRhlbJp7IQQ13+5XCyeXOQIMt6QNw07U56/tyTWzdETc/GfriSx79sO0
st45ifpzzyztmhVbsG0ztA/l7WvzCprQsw/2r3VbYKhFwaiFr9RbGUcvt0iXMxpR
PeExOm15466zEMlRHgnChLi1NspPacc7bjktM7SFZibJBYoXiIPUMYYQikq8THab
X+mOJpPFTQeXdbSjGFn4ESjr9EpDBafR45D/3+7fq4hmb8gEBngu+L6veKeNjPPx
LN2c/rY5tbpmYUtsnMryewia0+AmIoiyunz+/t7qpXITl2o2CZz0n6X2f+9/iE1M
RQ/tJoF6nHGwdRY9agWp2QAx8V0zgyZcLTO1RlZxOZUEvvFiiNAdGgs0uIupIDTc
1e11RaX7SmCNyrNvPc/qiBHiPOwQktJGoOWXleYzd3uA3QOGZy/3lmtEfgkcY4Fy
qey+K1I245HGNVqnejhpjyFVYV/3upg2oGTSihaNhmUFmLJvOgZ6EcR2LdZlRz4K
xlMhrgXHUyyQqESp066QAm4w9JG5tY7BqxrKHTzaCjSIc2QY6ZB7JAX5TIpdCw6n
MEvIrcSCi2LogBvF5MhYfckqLHdta4kBV8DHoYoRJWv1vvOD5rKiDEhjpSXa79C8
OiL3/JR7vhqRlLk4DdN9mdzqUvn9eWLuMGciftNQAO4c1bsq0HDluImnjSNNZTv/
Bchy4IkxqQ2FzYDpo+saadMZR6vNZHuG7hqXFVyrtwY9QMQVBWOlDP6q1JQPZXbd
gpXC4AyDBkpjt0+Ygbeyjly3Jlb6HQ+FP2aeNWWYYNpt+P0xX+zxbjGkDgjFs4Qi
8HPS7t3SN332K+Xonnz+GBvLlN5aoL94K9jIKr2quwA+ZxOH1OlJP5SNWRlT5mpJ
sB/d1ff75mDDaLxWLXuptzMj0TbiMj7C/hPsiJf9zOd0zZauhN9an7VYhhbhOtGU
eHiuDJoWlt552HOak12yotlCy4lMIrn7ux6T9mL3LVMZNvvjWZBRMf9crLGydLsu
3DxH4wpSr453XrxXzE3hHPT2kS3S83N3BmTe/joV63jX92kL8R714KAVnMANHnZZ
9E7poOMC4hDuNyRaB0pcimxZtAeupILX20W2Pkcbsrsi04fZMwblLgtm2Sa6k+SV
FLcxnOwYMipiKYhBb3EpXkHTkK3ufFp6VwEy21Nq67e3cJoIkLWD3Qeyi4Ozq6vp
1ppfCmTOHOysllKStKgT12Hs80J4vxi50qEkhrp/vqt5xoEwcHgqd4/RuDTaLkPE
pXeAmBfTWCoha8cy5Q9jZgBRxILYPTWSukR3GgckVcLB6YuAwqPzDKAkLLIUIQAG
vyg2cxjsS4jt3VnUI4HC7oN7B2QU7NfzKS17r/1VQWNuXQqKTI7hBgWLitPMwwN5
V7++Uq5XpzEO225scxxXJpWglVOeLmgMwvXac25OeAypLe3cq1AeCTy0br1YlSNF
Y4gvZaNwnlwBpmReAB3w5j4sSJ9JG6PKaltGXvU4WA24jsL7dkkAoFPkWj+sNGCr
jWpRa7tnP6JSZQb3WFAmgRWJue37BlbV7IPhMixVKldd6E/GV1xcGh3qfV72mN4K
Nt3MqJrnNW/Xhh9VAKsbcj+0GWiWNQeUlKe74XYB5MumLcT/W+p9d1PqhD8owKxb
ur+66T70wAd+aK3OxGG01gStcualBCUyhCSMjQFpTS869cNwc4VvUBN8iC+toO6h
dY38dyzbAPg21rF9eIY1MTUCtZlbm5P4dEa0BM2PEOvSHAuP8Yl0Q8QLz06I0zXC
duUl1Vau8TlXvWY2iLJmhEokJF+CSLNvkFUvJ4K9yvx+OAwuGUZJNBrBfalVru2E
CsGf6RV0Y/UmwyIr18T8WfemZUYv1S3iZsaCWKfS0l4IBgxaqxd0KlhXf+ZaLHpr
Z91lc+x2WXvHngphvvYBwfFHbCi5OtLJhYFzQM6dc3MdHZMYx/LbpLk50FJhdNNj
Y2Zwgljloc4JE349zOEyQJwLZc/AizsBpq5NeHgykUkSaF3LRrZtvuqNBk9yBpWs
k8ihxDSQPoSVDSxdmDBq99MbHHogHSXzPW7g7aYsAnQxgQJM7XCIqgIYWZxhJDV7
5kPDIWZ7vIFk6pV5YwDNN9mEfbLOK1Varm1WShvOnW/XaAPZujNBrW85bfg84F0O
1PdWOGpnbLYltS/41UpJE4thdY/zLfMQQKx26tFZ0vulI7LL9ExrF3oLzT2gNZCl
hVSQSGweEUbUxmhHjDEDZI8+BY9LKXtVl/iOInrmoDU3UDvcfbImuRU1rzJc70PZ
04asr82BvtH/8gw1FSN3pVcdsQsOP0A6L3I+6MiNBMYpcAnLt9Xa7jDSdjrcusDU
iRcxYeLTPQhPw+UvD0q516SAkmss7BZxxH8IQMOlPt3mRCEYGcELD1up4Ae9fmVc
3wEhozLgvx5mOHhpi/5YZUv5ytbFl3t4+pXCknZ7uV6fJ//K9hFQyP0eCRt1e2Xy
NTWnAkf5tD7LL8qg+yXodyggoTuKpAwU2kwgC1r5ZtWc0dUu/vPLIPCrQVQmUW8w
Vuia/PdqsB7ITmVPRYeTw29nmiuuQjbrVPKELyS02gJ+beEc03pH06IhDWOUvmhq
sClj2iKZkvkxpR/6d/AyZb3j/AATdcPJXuajKIHNTdUbp8hKOP0rzXvuz23EMSJr
U1OplLFGXpjMsHxqhSigOQJQVTydgJyEtEXeojuAUAaYLx3HhiIvygz0zQN73amt
CB/ahInFZq5YqwFZT6B8jcWV8oDv9ZBb+vYwDKrhnZVOZ09TVlPsSj5UW8DFUl/P
cPlFGyKZhb8jCCvMI1k6wn9WqFt3Bcut1iT0UnPpkUhymWM8q+74vTj0QYcXkk+k
9PR7E2xTuT7FsPbTE8YoL9dNgez9eZ7lUNj51KknPOSF2OhKjg40o3i1MgUbdrtn
yOsCny3YK8UtFAFXT//cgeJ7UiuEt8LcsC9zHaMSMtboEig8E+LdIz5goMLLOvoY
1j5Y0XCvhYVpZYH+DxufyYOz+o01T+Bc55c5Np690wx50tcVloEDyy2AReuM4Xwa
FrDL1LIhaM05+N9BAClCRG/jPrRY//aQq5DvIHYBUABiU2TiJRw9SCQrERbO96/t
ze1qfux3Viug+U2EeSKQIEjc8Gt4AoqHaIE2fwg7kpmzaCSHAmBpGGHM+qLgYHPC
XzYVvUHVDgeCxOLUNAsJk/LpDUsMCMbWGrGHojqaH2v+HGBeM3Gg7ml7veD9Hcy1
VuiZo0l81Rtrnnk6FaOrocRQI4Ya5HyAg5mCihINckVzD9dxjPuJDkhrg4H4yCA3
5K7aWiIRDVu+hdzhcXPuEFKZWUfTtNdjNX0yhaOlvTDQaGU4KrxLnyVajDwt8g/C
OHSrQ1KLscNylqZ7eLKeBwtpdHSCRGdxkf/AuBWlcezQhmKNhSM4PdHEBS/frgmD
A8UOLYc1dooUXe7orDoQLzGFVhFWehbDCwnoFwT6e0DIB1tEa36f5wlfASSXUKE5
alQIqAeIqu3JQisggxtOoaHP33pL3uFMEhAcLu3R/22C3ElJyQ8eO/s7ZESMBIBx
RTfDuIkS3FI1cXHekGR7lOIrCMITzqaQM/XuJJmU+ImTXKpIKtA2hU30gZGQjiJ6
8lIqk7kBxglLoqa9T8zRacMLqdhvUPKMQjAw9SVjtmw4/Lmb4RBS4M7NguH8Xr6t
SswlGMvR69Hyy52Zj8RZKAqy5OJMl54w6N38jgtEFKSUb3fq4418kdYS4imUVH17
+7LKNZW2Dog1DkowovSXVw/2e562UxV19oWIzoZwaRCQm2jEXte/b3mehqPTmz41
oSuhRwXLy8k5+Sm1Elebq8EuKkb8g16haGX2oWZJXQNo3eqfFJnhwuDmCNa+1BHH
3dcY+ne2szZXzREJNvFy+mFoBKk1oJdUhdwrlvfm91BPMru64uC0FvS/eL18LaFm
hseDNZvpI4zdALjd9HY2npi7VuyOtxDmbOLfWmX+VIKJi8U0+E2bITNcgaxWmTAZ
Sn38YHw/Njk3C48rTaMSXe0a2aehApZ+8e2Hh93qXVLiFslLPTbXKdoKA33lc1ub
O+UL1wopEK5kYxwi/yZvkpSwPkdQWrgaE5sZckWR5lPsXEP5gI/zy7bAFneKIiXl
n1enTFtYzCs10Qt0kUUOOi2cnnPgGEEfHPhxrltyubQapnd91TCKBSeTGQRuCZ6O
r6AQLwPJij13geA5PqlOgNPmUQP0Gr3xNDau1klDg6AqUuRPHYxEoF4BfTP8xoRu
LOcIpup4dFTeRG/oXTomtPGRSh7CuLH/g4KG8G6T+gf8M5FfIuyRB/pNWBxWRIxX
OnXHPjtEZNBzTn9rjRH6whLMXiBAwyd6MHbVO71hHeldUA8L73kLYLeB5DiZFRKj
hPSUxYtm3RqFfuh37nGr/dMpmIsItwHPzGA331yPXqdZgjBf44rPVu8emRmlBrS8
D1YKdzcRd5jAbL3r5xBC6F3watsE9NbTG+9pAbJ9vaTrRj9yzvCo0kiHU38hV2t1
ZLXtt9Ek4xj8hiWzmhd7JpV6vrtegLGOprpGaR1wOKYxDi7GHzKq9yqRemd3+q4P
IJd85eEuKP/fOd0UtaSogqjKPny7XuK6QMIthdCHcgOSWmLM+4OSpfGexqDwS+KI
vLghUKVUvu1MuHFuYW1Znpb7WuOzCgdTp5+YoZU34v6HPdMBnAL0Gyu07dZO1etQ
TPTcwVCWEfLrwDHlPeaIwv6+IPcs+Nmb2o08NBoOXaRyUeDFq+yUuEI7tUPiDRHK
Le2KSAaT8R3Hu4Sgn1w08M62CbJtdpng8VnTh0X+flYsdEKgSsaQegE3SQUqdPvs
WMiedzgiw/slZKoROLuuZVI7mD0tQtP4y6GTsiplLlwE9/2FGMGB+ldyRpreyTyf
/Dd3JXONqZqxRSjwulK0S5Sh0Lzmli/3049+roKUPTCnrEhQ5w/QGeb6G2Du+JOL
eXFOTdD/HEZ4kq1rkmB2rCtzw80XZATnGDIWXQG/P2c2e5sG95WqEH9L4QP72JFY
RFIOfk7tZ4v8Lf1PXWfSZpk6y6qezuAQ14Z4ptIi+EHhN0hvu2Du1sjnQiMaCO9M
3r9cEm0Yw4JVBgt3mQZMQya+NQza2wOV7+Cmh7B3GRXXTXVqTgs0HviUsCS82mQv
nt8yqo5fAB7wQxdM3325Bcm2Y1XKmTQWNZxLpLATGxm22w2Z/XRWdDr0kAqmyzDQ
zIu9tteklqANR+Sz3CN+ojNULpORldg251II1EQ10WF63sjDWsRHaJ+9oSzGG76/
3qrGhYbKF+O55ua57EmZ5Fkz1l7i/QCXqhCdvhE3eFFXxgWxxM3afiWh1aZePOG/
wdHVl99cHLNSUWQFCRCCpWfzBxJSIU6YeG0BGPiQhaITyAwGPVx4TCpjnFROAKWW
75TfB/HzxthhoVSxlC3bzNQPLJbltJ9S72AyLK1zY5JSNBTrvbXNloYbsxS63+pN
EGV1NA4P40k7QvoyCt0o51yMbVd+9vXYNtqbXF/AKgHZru1iSBack8LYHG+1izoG
lJNqrYeRxfI0oQD5TgK99MsGNMfWbGIY3bOPrelbr+gpr7zaNThEkeV1o+ZpGuJF
6xaMKw/B7RKC+kAaqj78hXaIjqt8MrAuZUqDznZF/PAZkP3YUP0LBEQdh7RrmLgk
NXhWiO7zn3CprKRiBbF1+q7VCiN79wwRy5Ny1CO/QWcQOsujK+9fqdLOVlT6055j
E/+uCNWj2jcJdsoISD3OmRBygwk6IMt39WzaZGFOU4MKM+hWHHwVlZS/rsxiIL+F
XCYKri0kFjtUNNLB7ecxFlqcEtyNDJbN2OrA7+qQJZOqpV4z31UuK7X893inQeNp
IhE/H5TKsC5zI7ABgFTnY+IzC+Rdd2892lc5wwrDW8Ug5UW9G0SKzighIcCBH5KU
hStlHv0PYUoAD3n4nVgUq9ncw457Bc7ezv9GmScrDla1G4hXNm+EV2X2l1+JXUlD
k3dnV2OpffhFBZPu1oLvC4/CO8ykP4vhIBjc7fZHW20hRWurcPcjj6zFwsCFWRN+
+ZI+g+/VNx0W4K4qewwrTI6fmWSsOZ0Q76HvYoaNVH26H9yjfJmHgDyoGxLUyXdx
DTbgAz0mpp7YSRNRGESY7ujRYl2QIZHyzWnFIDhhbUK+uIZ53FszEGtUNKDFJj+K
DfLvwubu4kFp6eF7hc1mGWslTT+7snJvoJG8AFDxiGx2JBQD6qFIlf9a4Hz17nb7
iWZZuhOsX3E1F6CsuRfL9h5r54EKJz+CptLkxIcqv+3KYTxV8z66n2J7ISUHkxoa
oQ3gw4XphTe1i71d0R+p/4BcAKdJLfw9tXAxkSjQzmIzYY6DadWRkj6lXTZPeK1i
1gyNh+TdclcebKLS2gdoTXGr3mRar0VXGGcPxGUo3GkA0e2D61rumC4LND476BqC
nxGekPttdt2x7z57P9FTwZyhyIZ+ZauWIWKa00PQyHn4rdRbI90gJRL3zn6qvAJl
gc18qniBM75wwB761UBDlbdwAlhohpnAODVQRrHAfs7gVWsxcYq4ndIp3/Wg3so5
ISvFCvN6trc00ZAs5QsRhc4BlW6dpdqeyCqw/zNYM+0HPkfltj6To2R7bzekAtrG
DWnplkH3BkI4iUQoSYcgp5ZC/lWNswcDWfALOOE9rIifXmTG16pQIWeLuxZMi9ul
8XYWUcXN9t/XUeQ2FfXC5LrQFCzu1hpkggS+4lYKXPoV1uTkpgcbBttf5rrbduB5
v3srXm+4Ys28TyBJlhkAdAli7Wjxl9kc7zDY6KhpsWVRK2bWk2x14ivPyjRsFL9I
tj5kSRxEa5XR2F8d6vsaSrO7nZBWf/56L+6oIFvaaPO8A9TRMnxiS3kCgbMjHfJF
NYITTFlME8qTE340AX0aR6k2XGcxBMyik2NY4k6r0GFSuxlJJhK7tzoj0YbmZcsj
tGTzztXgpaIDA1YRp9jCTXg6MiVJI05goppCYEdOIk1Rfu6PA+AFRTHl/FEJEQNf
F0F1Y55bcmaVgM7hPrjk6Ob497ACHLuYPRGWiTX1/d4YvXoVy87Xnk3TLCKmeabD
QsmieZ5lDX5Yy6WxPbtqdzJPlXcUIVO+U+ejfnD0dmaXqozIAjuA547rObUQQxVt
FApeMQE0oJS+aYZc0GnKFYjnnfvTQTNiISVnKBJcFwxSNvJkQC3j2TdkF4ACvuY5
KXnAYCSLLzS47BQElxmHE/xImjubSrXb67wc2+U73WLLuudp38i82hcyxG20dAIa
UtiQRitH6zMW6kMTNu8KkhtrptNXwwxyi22qzHluW0p4OaPuXrfF9QpjRz/3rGI2
OyCxhIooqd8lczzOjYpGebhLukx7frLJkdm4b2+wiRnnZakBMSfYDJsvJVKLF7Lw
eAQ76QNmVfjkFfvxeBLTdmIT6nE4Fbddsc2iUxnfSJ2V2f5chsfqTTtPSsoCMhrR
ozGVt1IHzB7+0PWJXmJoMbU0/4vfiTvyCLDhK4f5GlpIbcdh7w3LXpzU4qz4umZJ
fNBOJNfINgTUrfGHbohqyRbO440GkMlMwQYUOwR3eE2uRaF+0ySTlZqISqrMipwO
soYA3KUzIjIofLSF7uKrWEqkZxfe6240DsICSAQwXd8DteUUMpLiPdoJJ+MNkWyK
YxAnvmT6xUu1WrDPI+z9Nf1Fs0OnzTMPS/SgtTL7afowkO7HdfIEgKZZCbGt11hk
EWQmQyIZfJg/Wr0WLpjj/Ail6n04qaGxBqT8Attfiyfl/k4OzmubeOU5+jyjLnU3
FEni78d58rw2epUKZYH2ZCwi0DqPJS5BIe9Jh37JniMLZItqQ2wm8mAOqcIoU6yZ
OND4kphf54jh85Weqt8yq7IP4WMP8DDmwbFxaEfARgQvWGkIdcAkuRKRBHpdqKKJ
KcNasxBki2kSfFBxAoQTY3gpTnV0PbpevLLbDVT5P+Gd9jRDCuJY9LWgtbgbts5F
0yljAzrG81yQt3vLkmtlCfWT+GL5bBVxBdAOATSvUxktqhxUrcTnJHPK8ILxeK1u
h8843kRwakRlxrZvYG0KkPUFBrSTc6iXYf031W751BJfqCRP7K6GuezJjS56pAxi
NERG0vSOwDICKSw6hNUMkEDmnQIBtlNbdh0Pcy6jecF6mR2aAj4UkzOlStRvLPyn
j3rSMQBGVoz+Gjj0CMhwP1jfx0Yud0KiIlKboKI4+vvxU0PYpB6JA1jkq1ML3glU
6fgYDOkH06wwdEpwIxKoOfo01NwMlTX5sD7Wj13eSwgq3InMwDfn9eTs8t4wgFux
f7W5awvfZ/2t+B+da6Si5nK2EWpXIrhMu9rL1XCsuxW3uSRXBYfUcTvnwZnS4rDs
Fj+tZiZhALNeiiiqWk4vtsYnXfEyNaEzX/LNirBy3UASK6ziuD/Wv8yfgXNv6bnL
lvUl82Z4nHETAP54ALFJ7U8dUkFiYRkDXmGnbZpr9Rw9PG8F67od8SkpMmXsuXXN
XkXXg2525F5/HKb4uOHmsi0e/f12+Gy7BIsj2V8Zar5yGnvl5JjTCGmdxoTuMi8N
GQO0iG2t9CgDCSbsp5W+S6MrrOH4xurG8wILFx3PuPPIBuBDJhW4lccaDYKXmYcX
Iq/S7TVn+kykjCM3CYYF9tk8R6kqb4dVCN0b5QGCNOHtC13J0++gEUZwlGi5ss6D
vC2J7h9pNqjQwcYwCbcBpnV1MqFfnJrUKDHhqX56meI03DVjrZW4YVuIRFvLrfv7
hco63RWQuM0sdnDRziC2Qp7DLt4C3PeoYk8BTf3b1T5RTUdpfOGofZgczM6mRqxX
Ojc3QJb/y+3xVujMHxXmMpcs70ym1phuQ78rjAwvCMI6cyHqtPdIS3ugFmwr9e+j
a95YBQL+KscQZQt2WhqjYS9hgkHDFeHk8OWyIKWEUgoNONwzNYLRtJJpBumKCyg2
Wq2bno0nizdVra2AkNARDHXQJwwak/sspj/H99lfuudCIGyCBa/Tai1KIPZ8vXgL
q6TLG21H3zxn41OsqwgCk7h51/5vYVhPZj4dXg2MZMnAq9Ksxq0soMDGaQ/e4ezM
lh1vt4tA6F5wnhT8Nm5gmkatHvw4//h48psB2qQHLuIpr1Z/VD1hqrkqle6eKF9b
sONRZnrzQ3s/m8ElCcN8Qjwk0PeMeCWRWz3/oLwypdA9vPYjiKk/cpvR2+eAQvTC
unqF3keH77YTzLpIOZW3ml2NEcsHyXI2MMc+5/XRgq423TpzQnYEr52WZ0hf36RK
Zu1keuM6khbgNf0iUjm6x8OZEM1o9xU7sU74KHHaHy3E6ogmps8Xq5EuhwZeHuMh
ThVYlltMZdoeCvqE11f3KoWqgo4nEuPyLFrzXDkryymIsumS7GLehvVt+DEqcVCG
QuOyzpzoWAiPfqwqrRBIrctcsTsArfAbtIdT5g6AxOuhQzuG6y0XaCFiO/OvMBdJ
WOaEGvpCShpOdBWB3jgM5V3kzSmMUStUOVqaPiL6as0nYb7jcFyvvWyR5OWTsAt+
Y264GxxXUCPhtItT6xPl+vwZzpwcXIiyaPppOqBqo1e6KYoko3wzMQOUqsIqCWLz
gsesmkG7atjQIztAbNyw6ZRBV1A//D5pPc2cYLAKWfEY9XgKAozoLfVPbXfST4Xk
J/GGgw8O6sBmuCnrw2p04GIdvnQQB0DcJPWpO2PcyJH074dvZYgiz9OECYCXsSsK
DRSYB3P4LHnkD2ap78e3Zj8Ywx55I4guN1tNcXVpjXeakxA5iMW11OmtnnWkHgzH
w+IOFX6uiJUp5PuwUq66MuR+c0G6VotExKK7fifxVFE0n5MwPb8Z06RuOJ3E5ghQ
yf/zsNO0GJJRDJttbFMZ7vlPI9Ckxs3XQYItfaqRdU4Xn4VgtqFhDJUEG3cHMhqY
2xSkoJk+bQ9g1yTMYcstbF2EIdqo+DUxdpyhn/KXOSVH4MZ6/uJDh8QAWWmOtBcI
bmhW7kIomJbFvRGwwyxaLbOOpuHYYvyIq53+iGxTtaGWnHiOOWn/7s89XVBrqE+r
nbAHNEKMHI5C3msIz2ltoE/LpnvHhdbR+KYAZSEru+ZaKCaGILXmwFi/7hDHJdqX
noQ1agJ/cNBf0938MJVmJhrY8Z3TJcc9UWSuggftPpT8sNlSc+pxblbaq/em3HdC
w0nfIS6mE1n+OOSIRPRfpfiVY03oucu4P5ghfPEjxKE2g3SsnOr10U4maY68wp9O
Smk4hAlwUQaCUX4y4SCjljTnI7U0CIH2RXDx+hf1uGbx484CyIsWurITTf1A9yki
fruiYsZMkRv8pf7L6CfxW/0mVMTme93Ungxj+Wm20G9j+3hQ77EHgafjikEgd5lh
OhTAotccnPfk1mNAXeOnkcaVhGpLE1M9RQlL3+2G2hY1tPo5pTpDy6mR3f4KIWxo
FAj8o92qXs5ViM5BZjae8ZOC7nCOfRkE5G1awKCyEtmkSYHJkK6ryXmFf45XbZOp
prJQPvU+VGhsp5jD+ObNfmTLPHvGgCJi8zOIN8TunVX7by4/UJE4s64ePNhJYsYC
T+xpicuL2AQGf3Zwh4Uac2hqeNEYSUaik7EC97JuoBWIsnUeSOS0l2wmviXIq3fN
xf7Umd55abhNls982uaI95IgKuDVnzXqyt55pMOBK+0qoWzwP524kr/iNj6YLjrM
W7K3TXVKjPQ8ReEJLUFbYBaWWtLU1NHB8epegsPzmE8+Ts+e7eylL8byEUgnY2Xl
Ng8bm/u2VnYsQhHlMMim+Z02ESiI5UnrICTTFFwxsEx1d5z0BHm9q5MBP5Mq2Ug9
Wg5i+eyZDBVXbqA+di0DR5fEBnxcDu5tfYR/1RN4fBvTzGC+njGBKEb7EZ5xeftn
zMHLkB/gcfVEkBqEvJg+so8oYMEGe2uP3pbcWfju5tww4nDOfX+RiGqAvmGZ7gQ9
B+T0EIkARIFwc6UafqDmUQ1x8CAv6uooe3mkGCUSXsS1m33Kpp5YOiubsASXNA12
WYZDkqyNhR7JHW/dIJbiPkF9ffR5Mho20BbhDoHB9sypZ4qsUgUfn//3PnaoW9xT
sDrTUtfliQowAOZCH2ToiH2pFS2UDmU4VDuqqYI5ZAReNbfELq7758Ifu0ZLwvcG
RDhblsUONlvujklx9CWGNNt0VwHUmXGWMmXYd0xDaxh/fJKZlVsfqj+oTgHc7s9u
ZnLZv85LrXyWlmSfWKbmFJMDg9bkOiqP5OLqLvlKWwEbcpzoEqEuGU+KcTsaKBkH
woK7R6JtUt8qW3OKFI1FIz9+1gtNv9bBeaFFaEtDYEHgXM5Zxaitxb/YmB8enuYk
XivQQGYXzsBODkbWhsSFzx4CguTqK6EKyXFb5IiMHZRK/FadgaA3VJQ0wTd1deWv
ENTbHrYg5XLWaRwV8CRFERBWW0j/GUP92miq4DaCp9n37QKOcDtZFtzAgvVbDxJo
abe2B7x4PsTrB2xDqkSCXTDejCPS6vW+IjkzX8xzzeNq65oED3ZoqcU092qOmUHF
mjymqEQv6y/09PBJVRdebYyPipS+FYjGH02/U+OUGRQTtye7vPgdX12J6VwEsbvE
20BxLQ8ItNxqyH5RNeclWNOE1lECHAY88D6ytvO79fA/AjttE6JnnGloU9VSwJ3u
/j7b4Rf5mAJybrQ17HZmGdXLdjz6N+GMDJ+M8T8L0N9k4qZ/l4AbYFCqJrAbREsS
1wRgZJ3lnSJKbdH2FOnDBqj+VANg+qxBE9fPaSEJjWgz8ttP0pJdQZQW+giy5bd/
hC7NSPmzvye10NtcyUGgKKIk91i95n/OOAvVKDYYUbZ6faqBDYgMMvhR1NHselfV
/p6oEQWovjC/0UUHxUti/uTILYQ+Kbvf8rNAJ/KH9bBqZQPzZBLmuK81NJwZMt1T
lvzplm0HCVhf+6HAVqcob+V/aO8SJQhoG/eHkzru9gFeltpHMQ2RztbxlT7fDyH5
GyE/803cc6SfclYVRLJtJop/qtIqci8JBc1OXhAPTWTPTwuq2kRHuj8uJNeML+nC
eXi0+0Tq9mDi01DFhuO637LTz2GCNduG02ATdNi8eCH2esVmjBiffZ2Gst5AJxIL
2R3cJqyB+B7YvwFTEWX/nRFBRXuEZ2fFfdATWAYvqzHWtxEnz1nrs7BiJjkKyH3v
UIdyssVsseMtAgpndm6f1BMf0MMuDwBfYG3ZD8G+jIEwLKpF0kps6MuQEExUyPYA
JM3xq8KK7HjwlmtdAqkDpiDmga0cW2KfMfsKfFxqJsz/nV0rOQqimctRhjPTgmsT
Js3zj6yanXN4pUBkChgGRUB8I3uUL229vYLoLFk9eH8g528xcSXUJRXzCGz7N+bV
QWCWKXvfxVVfb59GmJaRD0Y+eAOyCcPY4Mc4vHaC+Hc3rcNvpCRZGVjy89kh6Yic
1SFD7LamjDP06zt/UB1B2y/JwsaWa23IPPoricfIT5XaZMlUwr8IpYRGibgLQmvt
OOxrMI2otYWJJcZ+Lm/UQZy8BUm/n/O2D+cmAAssc1tN3LyeleALoKma1jrIbbtf
y6+SRg/pyR1lnU9hcKVUbc6U1PwD5/pUmD8aGaD8LyZoQDsZ9ir7GWW3mfz27Ugn
eUfDU16+w8vz1AYvaY1EbyjEzP1GPTnVEGb6fZbXTwJeyk3ilmDfALJ9qvdLuzsz
tlykbml352YecpRUd98GsVlocrOB/QVdbeeSPfAiHpp5UhUCxSoAfwGFVI749Xka
CZ5+Djjv8O32+43tuY3uT+4ZQe+ZnpJxaK9m/6XmWg9Eq1SMiLaOexoffVSoIp87
/5RlbAI3Xo8j2xOLbs9h6aIBAPFR6g79DnNj02A+N/gZESJOU2FvDaDexapcFDSI
lj9a0gpGY/oSnEte8oG7QLeYY19NsUhqu3UkFitKTFz9oXnrQxPVjW9c6hBpTlbl
SIv2yLwcr0kKOL3nkvGZ6P67xTiaU5eyb7izec4dwvhLhmB6TMTDv1mJ2sEzc7HY
duKhoAQpV9UqKhK3Vd+8fV0cNvtKWu8unctzjeCuFqrPDEbtg7XVWgkr0BfU+KEQ
jZ6WEedv2xBnURKxlJHfIo3pluSWzHcddfe1aRCJEE94EyZ/Mf1XEZNFc1JJIzd4
yG9FPKN/EYn8fm+hGOWSpFBgHCoiW5QJeGB4ba4HKk8W71ULOJ0WE4FJ+HxQuXJx
4QEadR9ZQdnVoK0VlSUArqvN/Bxg+ehOWI7THWPP5NNNl774aq2ua/mnlvtWvGDG
YFKCuQa2DSkh3V+IrY2ndSPmUXTZrQBOebfcPVqWTkgscswfo14n0WK2a/mj1f3v
P491tqPFc6NOQMwRCnbnRCoZAiSjCtC3k4Mjwp3fKnwTavhvyy2Z+6NReDS5uOwh
XO6lsmuU16WoGEIMPcaDcPeboTlT9rfLz0Li/s1qIhbs3Ch2QhmyAle+uMs7a1ro
QNB77ujv9KCw/UsWMC+KtVyugjNyVWWiuBKTmqu6mpiUJPK6RlzH073Bo4FJsttX
VYJWsoknhuvsaUu/BfWKkoVCkfGatyavoWPV8Z69AkRjzsUUJzKkPwCWUFV/fGuG
vGhQ9Q+D9CmIR+88aGcCSPVgJye54w/S1J4aRZZ9ij2GkePSqiTwiYmqEwgnktOG
QfPdbAKw2LY4I62mJD1h8xc/xTYvLlq6fr/4HqjdYeNJY9y5oHXI0VQZOCJXgbAV
2Ny3nohkRCqW4pWli66NUbzg9ZhW517iF7320nENKdtM34mE+z7ozBTFFLTCmVqu
QO+RkReiMfHIkPQZAA2sP+UeP/VRk4xW2WCTKHSOQ4ayxneTYk2DVdI/lFQ93Kzk
1T68p9a+uw7NbWkIr0pOKeEf7ysXwhmxXlkFZF4/iprdEcsE7Uwvoxy4faaygP9n
kmYt53xib6zF32mWnPX9AbQnVNIxLNHl+z/28RlS9Ia+nKCWx0SWGtkuzl4jUSSH
bB1hklU++F3CoVTrpz3l75x4sGSCe+HEF8YRBb/zmYObu5lTXskakgcdRwxkTU+h
tdKA6yVRink6SKlTGmATswu22aQD8m7l1u/jcquXmc4d22P/vQzN2Lg6bjVAqD/c
4+n9MKDsyzrmjGrASl1obdEFmLH0xoN4buTdC2i4OHKch8PjmYoy2oV74QCytwJL
hJyYsl3Wjwm0UJ5TALR0OaVXc00RE+EVMwXuEbROtRzC3MGr7HALv7yqhpKf7e7B
Tx9iKtFRC+C+lV23sRJvVy5T4nEN02vUm7F5yeyM6uiYgGMVljrIBqpxKthbo43f
V0NQaH3YFUPv6gHO3X1QxN6KGqKlgs6i6ODrP5o2VeCKFRvElbT6xf5aGy9NSNG/
Hk/th61Zn5AUFB/aumrLEI1GvlgNC90hys791hj5iIo5dyytTtonwjpgkvFsMo8B
6kFpSq6WUVRSdzX1fVYFRkwWy47M5VnZOx7Lrw4oO5f3dloBwfBGPv143JkXFOcW
G/XfzKHZxGHnR/EXGbJgdyWlbinMFpuL8PlaZ9ZB7EdgTYUPcpDJL6eRI9p0nP02
YZNV/y1dunB6foyd8vtaVM9KjxiVjXVCZtjDadGPqvhuyEDPxnmVrXKd3asUTc8s
TxFVU7dDlWePA2PVBpM8sCW4ryi1ZaGZHib1PTFWWU2Fzm5RN2YMxvn9vN8YabyI
u/uH2rqMnWDFfC7L0XgNNY6DChG5+OLS6nT8by1r/v8iTl3ioLdw4Gt29kuXaUoc
wNoUySYOPyxNZNlgoF8WIl5A7pJk8qp+BMfSrRY25FDua5pZjkBgn75nG2wMKABP
uA8lnA3QbdQXRu6uE4kYHSf4UR+o2DCObEYt78TuKjV2kLVu5qUly6gLoIoo+zFK
JflxxurxUJNxsHtsrtrwhSSPwGT1icKe6lyiFgy28el9BN9YoJbJ2aCQnTp7pGK+
WPZlxSP+c49eAFgsEwC5aQu/9oYLhlCl9PToH2Gl/We7eE5sjdYAVxZMysPvcbgW
1xKUTXatJlqfLezSaeJ1XLkpAENUSo99l2yIZ2tTIM+qqjdaaitGUhOSRcn/VLt3
qkIhbTFsn8A0A5FMNMgX1JHGXNHMWtfpTbKrktwATZP5rpyl2cRBK7Wr/9JA/KHB
e2VbwixYjU0aeOlG3ZwDPXeMcpeQo3Nrg37WVpzc/VbuusYis8iuOlttRyVYyE/a
62f+3XtprIBheTaGshB3uUZwj2H4lh2PyBRPyJDANtlhtlqkKNRcIjDLILHDwo6y
K3zL9ASwVfA6AkgiBEJp+6ZpTEFSuaNYrZ+J8JJasIAasrqDuOfIvtF8yq7eF0OV
dtlH82JW3XMAfakc/aNoK3GvvtYk9A0Yf0n4cTBm7w4DdUXt/g6Yd/SlYXtfRWHo
c8qUCGiZNfjyced0jIKzCvC0wD8b9rcPh4VVGWkg+5JJL9HaNnhQyTtgVYcTc7lS
7lipyVtLfDlPtNvl1bB0E8kDER9lZAmwurXB0NoFiGJ6W32kkWYWmFofpXD4dRjb
0PgztArnm3qigZ1o1itCVF8OFgLmfA6g8MWYMQAVQsOXGj0wTa6yy1BIsmKbNqsJ
UH1Kk18LaXC3/KXMnq+QhA3+gegGV+/AqsZ12yENM93DkcoPEuwJbmlE9lr2CNfb
wm33+OckKVTvhfednNwoKOAEWGDtywxw/H+BWTGRT4F6kYEjxhv1jnQUGIQFmf24
l+DqBnLgtlM4gfha0jqQ8YL/FLck7MGsXWXV0iNXeqH844S4LzMnTVgJcoddUGKI
z9enKME7+wUhKlAP7B401lpC8SMxIGKGp8TxsFN9s1RVdG+tUrkBQq1OBqcsgzlU
7Pz4k3AOaGVH/CGZJe9YssMep4sa7A9rbJrbOC8FckZKJzNsQ6Fticrg7yyjcZ8G
D9hRKtWk/UXbxQT2ItL1r8OE3yJxI+O8FTo+mi5lfYvyMc7htdsonWX6CU6DRYoe
JF9onSgg3x+mSwv5yzLO/IzZDpQ1G84qYbykuLoPOhU+oGOpjSgNZF63Jef7c4f4
rSivNGh/iPXwt0u/xbFV4CbCNH+J6/CyWmJshWH4+dAnIDtovxE2gSCtxbEWq+rd
Ynu4EW8uu0/KqmO9fCJ43ONYRzlDxp0Dh40D2qQWKL6Oldbl+kcqwqx4uKWugURw
H915NsU/pVSJkZq5GlZI4Gmsv85faLlXDGHoiyy2gHuC1kSfl9/+hTb5kVIK2VmR
xKetM16XRTNMow9tCr6yvTjLDbJ7lKnb/YoH+gPbWJlCJEcotNMe3UCQrsL7DvWu
q/sh6SXkE6eUZI85i2zEQRRkUxLZd7GycrkxPY641/1e/lX9jlUNFLtEcjsvtXbO
0c/2E1hCa422kMPzuL08iWibYq3LW6T1NTyg5uacnQi9MxWfCPc4oern9z9Hbazq
eExiWuAcSKzQxjGugOxEFpyfrlmoaReUomeuEdt52XvR3GegWhGRz4sfRG0waoQm
pRGb/X3WrzN4XHqSqnlEF1ksrv9/waaza68tM+dOCS8juFzdV2ykFYLkNZqgpvi8
cRARUIMPUiKvYYaXb5Q0XSNMG3l8K4uxzvPqYy4TNEIjWlmRKzpMGGSa2BLo0u71
WJyVWrggtwh1gAxH2eoRuQdCdZfWRmcPF7VcsAAWM2DPfo41u+NTOuE4UfgoWaqQ
Mv/vcedQrkOlUQimUNdRJYMURY4uaruYW5C+7jd45oPl/cnx72yy5OjwkdeJE5aB
dFS4NfBNtvNHYr4ZDzx+YsKRaxmzyxjn+pVg2A9Yyz5j0I8umfOCG/ym3Z3OXIea
36r/wT8lQ7MfWjp/GOegJwhM3JXDwj3H7s9hc3zmU1v1YNiuHX4gbcl6MVJCDqp+
Hm1kPmvxCzS8YN7Cx/CpsB/C5a4uHdmTo6PpvZBTzpraHyQ1I8xaXLghBpH9u6AH
bKT/BYAC4tfZ+Y1M2CuitmfESauJMrOA0d0ho3YkglV6hIx2l3/XA+Vx2Lwsswg0
ml+r8ryyryCtTcL92KB6IoZ5/xDJ7UuzGh0ZQ4ChuQzYMVa7aa7dHwEJwq265lQ0
2fCyjBV9GEKpmPrHTv+84ftO97jWQfMjYGEFlBy5WZRkBNOgovGFKggffB6uRNdC
cLjJB76hmkDz3HISIKr6bOdgqWh/dRPLVAX6cjRM8RrHFX1wD/D6DHxEjGDh5BWX
1lpgSgiIuuU1W3y5Bh43k8rGFnBxp6oHrxjDtSWeE9ZqCsqO1C9qaDDDF+qU+nqz
rL6/1p3hTyaH1GG+txgurAWJGnov9fYkvM84yjTBHn7U70h+DFINQtBP9oKz4otN
FJhA7qSJxFJQ0aGtXC14uiQY7NeM20PL+MhCBYsDH4bRlTnWy0OUVEqdSNLVoA1c
9/8KVBpAXrykK4fgRu4GWZBmhJh2ma0wzAFFQUEPavkoDfgp01gbzXhKLWvs/mai
KA7eE73J9L+AzSzWmzIhO4OZ4NrCrvzmU3DlbUHoPDby5epQy7VTxyHoQPnY9E4Q
3G+aolPVbAzBhp15u4Lmn3NMXVV6BrYoWNw2/4bH0vXyvInAhoanTUHWX19s6mH3
4XSft9xYF/88mx3okWn7jiHZxODP4M+57t33zHMusp5WrSMEoMfQlzcnXCDu9pxI
55TUuxt85hrSz4Idxeac6h8zGD26wf3xxJYBzz+wcuB3tgI81vPv09mviabv1aD6
NMrDFf/LAkz+DkUil39c+KvgJqHqJ3URsvk5bmJZlhO1HG8Mkrq9HbSI7lCdFElm
ew+rWWwpkQi7NcZnnia8cqtrmPRmC66R2bP3mfVlguhmqa67Z+/xMZAy6LhlOeU4
Nl165d/gLdyHr7+fezaE+MZ4pH1Q90N1nKK6vBU4N2+Gy1nwko1haoKxLAVtebo3
HYQoDwjQ/X3tghC+tOPP+DfB1tssPaPsTDoSE7CCgwlJP09PmWg9oRMqQRhl7igu
eiGPwzAxGIrRqDYTjEBu72Zk+zmi4t7HXO7wQo10Pxsgrn24TmYX9yyk5v8fK4fH
7I6SW2wEhxl3aODQbxNLMlkNjSQRjRA4B1PMG7lCK80gvombAezHNQNXfzra8p/S
999DuRB/3sik/mmPPEbKo8+S1ZfvV+d72o300r3X1eDwOBuLoqz+Q3Zfwmlf5NED
kDFTtMwORXPgseRJMESZVLQwCA2El0aDvgYC+aovB66P8ypXcgvRBDp6dnaadJk+
7bm3/xfojcWZFpU+WrQkUHyM8AD9HolG62OIwe+sndBjjk+C7DXkPPc9CPv2XeqW
IArJ3G3KqkTgx3RXxhNcrrBXnxYOD/5Lfmh8fxaBc78l9KVGOpqP4daqMAv8cYR6
31lSwye/h6jkjdW+ZYga14Nc9e3DElG8ny3JM31Qa5xfixT3dSKBb8xRN9OGzGHw
eQheYpHC/E7NlbGIUTs1c5NIeteUvNbFDmoElPuZ6u2o9CmkbFrPfStTNRLGFKpm
oGONRAlw3iHjcHVZ7C4bAc3GZS7bd/RooQQ8KjPfAQh9goP48B26vhG6jltpcNOo
qA6EMu2aPZTPL6S5PABVAgV6a4m4lpHbVWPLsolq7lQ0eCQeTFb5c5727NSyd08v
1au/VBoydCqQc7i5h+GreJoJmrYaW+C412VsndWuWjAHby3qoF2D78jsQHHiLzEC
fjoVzsGbZMenlmmrpCNiobmn26FAuMMlNKJvoCuT9RO+jDl7EGvRJZUeNyRglWVr
hS0Zp06Gq0k5s8ITOz8a/DNH5NnjWLaZUG07rUWmIzdXUrEkOXVGk3hkITEOz4DZ
ZFHXGZJrlg/a/hQCLOZDnsMAvsaSYWiU8Ik8N/bvDnLwH151a4VKrtPNOaHo3yEr
e24VSAXmoREfksh0SitTAutPq3zPFCGh1R46drsnq0SxELWn3gWeAC+AHcw756GW
J1c3vibK0AV7W7elJg3ZDNktZGQyLFnGjXUvXGLzmZkJgXIdimIAuwk1ZzypQJj9
HvFqD2oHcJmR+GG7pk2BUxYjUXZ2XrbcYVx2qIVO2KieTJsVUjqBqeP1UsfUUpM7
btO5dnTIbN71dtQXzsLqs66Nd92y6jiW3cX6shVS9vjAULx52bDtT2HEBBYsFJxR
wKp9Lee6HyermgLVjaM471bGJLPj9tlJIazTuWYRyvqKaw87cFa54m2s+pATBRH3
2HVgqy3WiEhnjLLqXikD6Roeo4JlfE9zEXogDceoIgzTks5gFJr8Vcp2TzaUsc78
hJam3CHk1H84jm+QOZukaG1VgvjFee5Hm+ue28D0iw08Ns7mRjU71pTCReqSxnOh
R931k9Y7JanYOsXxlCnr5b84Ae8LjXt7hhoFPCn2dfOCfVpC75W3PLXRCSVsAU8b
Dn0+JOf2THceKSZWgOYt6dAZP3iWrehc2wDObXu00MvaXu66qd6I4YLlc2z+IuFI
hMBLud1JemZJgmpOW9+F2I0nAgZw9xV5s3Xy6XS6e5pHa8km7jmJakhmVV7hftqa
MNk+PiEigobJBvA2XLvdmU5iIYwT/8riLr5pyLavXdPJb0VaXNVBq6ugkfLHDYgP
idS0lMui22sH7VMSODRx5bXlIssdMRAdE7WsTrY3WzMIMUuYSr2Ew++ysgvXAWIJ
qkIy46bgvtgXuMcQu5Yt4SXHfl6ZuVnFZ+6OkDGipi7d/dzqTsM3/R+aJVL6S25c
JEorqOaDtBZL1zZHcgwvvIGbmQ8MGGN2dSHIZnXYF1wIlPGATQjC8O8DDJLnYd84
+isSuwbMtXsaCHE3v+LnnLruEo2qzBfH6mI+QNwKWKz4TcMdgtXw5stp63nsttJK
WqKmAn5NcqYQADab5HIeclkEflpW/XVoB5P32xrGZwg1ctJitvUKp17aKc/M1r6f
kzw/4ZHj06vx+Zp4s5XzCkZpn5XjwmWmLXC+vJO6mIsxY5Cny02TpJkfW/ZXE1hJ
J3aJzMMech6eEf5IervKJfUOTLBY3179V928fTLquyJkVHSDWBmRoIIWF97luMTV
nbKq5kJFLxyGb+PtBJVzjXDzAsQ6UtnIX74IXST3tRK9Lnnf88YP8e32zu4McmVl
TYNT7y+yQuLwlxABdf7ePypzdz4zybLLXaTlfrPwvm6sajuqJuM81FrrTGOZXGe/
P1IvjuL5P4oSktfXOxiDVEjzXtJgF84o3uVqG+Zo2guLlkXwA1qsUjdWE6bQ/z86
9H+dzaHjqY1LgFyyawKXMmZXfdbMZsbepSAU4gFO85U0eGODAxdLg9QX9hbv1IJz
3VSZeUtFp5gjoTovq5wxqyizR2SxMI3+D3AllVcQHIpOTAiibNxIbOGx5zrJcLG3
iXDiqW6ArxdZCTnWXScrRDaxa6msM+0EPlM2+M19x4dBle8OD9Fk4nE419Z/OfYI
speQv3DziwmgnpO9RwuIK4taB7GCwWUljzPAs9zpMwZnKgbssr126ZhlLI1qUVG8
fBMCKVU6u1WHn7N4myvtP9JFc4g8knNW6Zo4EHPqaMPvZNk7erP631tOY+6WOa8Z
NGufPcSuK0bnXck4uwWkANH4JLTamfExa3ThwRkCuTPjoIPug9u2GLCkU78tvpfi
dmruzynMT1KQDvKq67aITz63kXyVCpPHimxs0fznKxeAQLOGKKUHkelSEHQ8a2vC
6949Ln1Xy+PkBbRafjWLRNKvv78FnsooTIHXVxhH088qpiQ+Dn+iIoQRn8o+0l3U
/nBBkKLq6HKlwJsg4nrCp89qztdqHcKXkj3MHlNwVmE=
`protect end_protected
