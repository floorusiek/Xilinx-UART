`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "W-2024.09-SP1 -- Dec 03, 2024"
`protect key_keyowner = "Xilinx"
`protect key_keyname = "xilinxt_2023_11"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
J9hOG7VfMLL6wnUPNmB9thWwCRRRisPsAX7O32BnJpn494Jh3zgwPr/C9qV3KoHu
WtjGYlQMIdqYD3N5NTkvKlBwjNpCeO+2n2Na84qsvt9KXybGvs09H8i60QyVWrMX
ftGi+Wfg0JrULWW7RwA7b8uOxuV7l0JKO3wK0mPVWWeio6FPDZ2TUO8hWktwtaLx
yRrVUaJ/vsuIw1lRORRwmi7a4d9qebpVVbqMtBaRd2q2uUIGaMAheDEqPEJof8aZ
4Yj6F8YhaMFJZVbasl+ZQh6IKn7CfLIcPHKqwotPLwRu4zYG3u68QsBXLLMjtrbP
rPC4F00HhBs8dTtbsH33+w==
`protect key_keyowner = "Siemens"
`protect key_keyname = "SIEMENS-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
Gdb/D70kh3mgSiaCNMg21LXvpfjllsYKBPBb8aiujfh1NWlK6Tt6pw/SrNJemtL6
Q5XBAPw2SqkjWZLr8BeoaFga8vNiT++M0pYHU9ykHjJ376l7+SZupcsqLnAYQg9R
NKIBEXUSLlTvfW0BdJA8psmMm1JfGheRwUagezc/s2kRJSv564VfsygKzsIj8Ug/
OUQSF9W8lDqonP434gINmMRSM5iuReCaYfUIrrlAuoqPg7KCKeTafOcSiIOlDM2E
pO5udzAL+a7QFwaK611lLP7o2psgs7niJNS314LanCNJadsMc/LLCj8slhnkOGcv
RNVkSVabN8stgWF4sBICaA==
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
fS/pcc/KAyjWXgPjGH9cHoxG4Gu2YBkWQulMQz+2Xsx/gMcY54iH9Agxtr9gnqLg
dMLP8y3Px6EzTp0jjVEwb/TtZy2hdQhEmbCIcrN7Zr4QF4HIYG+uT+lObDc7BPaF
UPFHwRzXlxJcbgNz/QB+BCdpr2Bwg/A+SZLClIpqa2c=
`protect data_method = "aes256-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 3728)
`protect data_block
inQHJWbkfBcUkY/YwzCfV2J4bFLyoGRLJWXstVJhMT8phJpfITys/2gmrW3OLZ31
3u0ZXwS6iEZ6lZmw0U6qwrAynp6ThoWTyOA90zpTpLX3SinZGVwTqtjCMqXTZrJl
3SiD/4HbOO0eqncU4vSNlcnCmslr3/XjXMzS1HXIoa/c24+muYpjgOxaEvOpTWZi
tpLcc65D7EjiG52gyFQGIYQueEILQt6oKx4bNUcWbjiXdszTKqpt12OpL4GVAWs5
bAr6WMA7wE80U+xo/ntHQVjhdt+g0/5f7mqGfYaD+jlwBtO13ykYjxhJ922989Uj
jqc5a4xzM7NjLAP97OZwG/YDCaQaJ3apimHanMu6hhAIiglaF43L1w7d2cY38vS1
aBbbJDFFHEar6BnmFl+3M3YGkMxfpOcV8L+6nqeiYmaf766ESEn1CG278eoW9NkQ
fKbrW6XbjYYjE9/HBG0ONZ794lP/bUuHanHv0F1TYUZX7PbOfx0MREp6/cFsFk6c
PKWVLcYJE+f661/GyDjnW0OFfyIwnj97AQ4i4rXGMkjKKcV+EuF2BiWNfwlTQnIl
1ReoBeAnBOlu93ozdtOGc+Bz/jXx1uWrSR8NY5YeQxUAGdNB3O98VM9UNAb1lTbr
IR4ZsLkzr+vgufQkS2JPNAG5E8rag/JMCtK+TnXUUlCrkudIPFqclJH2CQnhTK5B
TCXcrbNc3xABPVEVTikrL+gEOlghDIQm2EGzz3J7EcK5RvJflaK7pP85l735tOCB
3NAZtraTvdSYxyy4KjMRSHiRXisg2TCSY/C9kFrregUU/HMS6YlHk+c2sfySrl1l
Zp18pJKL8MQfpodvuMrgF9/bvK9ogiVj8cW0ej9OaEaOXzA3SBB5jaR/zmAciOx/
NZk/cURZkdgxZLDdrEt3ZBCNPzt3ZirIRYIEnZVkSMRLoHdgejEFJDd4SsQOwsED
zru4hBkNsVukSQY2GEbniqZ68HH2Da+vvzPQD9wpKFbpN/PcvzWA/yMNZ55xyX/+
1we1hxdfTiWLr9S+PMMvTvo2D0kIk8D8J6+nvDLeUy3/3VvflQTFJuu9ppmDe/Ab
x8F5q2/o36U3qJwXxzdGpUN1drEdQcILw/fsTp/Iqy+zBss6NwUhF/lWqxQPqR1J
JmtWLeaOYR6mlz7exkF595VCpu7f+MQzc32wVWOhC8A5u0AuvyRCFVEUAg90NakN
HtDMyzjkNONxPJonQpk8WdcFCNICujd6DvM2uEJf9A2d4MK+eQGaR9oiepOPvahZ
ULsMuARNvpqMHBua3EdBKygSUcPUFXaEWUtlZ9AtOQkcw6laoD0IIXJNovmOttTn
hCN86xTwAVVOrjfDG6D/GcT2oNAn2WWcgR9+VI5Yz6YGrTrccHD6ORc9289SB836
jVfH78Oj60f00PKw2ei22mp8iIW7Q0GptvBWM83TqvQgDEQhyhDuTu1TYI4wza2d
rZZaGpI/FiZEXA3AneaUgdOwnyq955h2MnzRvfRSfYxoZf4KukiXYQwpwBgbmecy
sb0R1Je4hfiTif0YE82cX80Rm+14BNWYBfFQATbFusTR89Zis3S9XVSkw08g8Hix
QJh6+Vs4fKqaW8R8/Vtvt0nF4NbO5Shp/OQWqVlU6QhDChJv/rh91UXR74PuiCgC
FhhLwv/bzl4b1yyUmHbApJ2drpl7JNfWL2UFDeXTXyFA+uT4a2HyDGj6kPJPZoD+
wMeI4Ldbtp8hNfNKO69CyTGUv93o2f+snuUYLIBFpLSPtf9E623N9VUyf2fdtfM7
tFG+wrUsv8XA4boljO6/ex/LKNtS39F//TO/X1afPMyOfhiUvgjVK9D4lun6OkcR
GxwKXrbVhsU41cftiAcgySquXxiu99yeoMvD0dmMvmTgyuvPqLpt8IyqQGLYTzK2
fisZu/fTCKUwsrnnuHf0vcBuh6ONqt2o8yM7bbHGcaJdZD/94CrW7+6J1bcOGiVt
TKL8ubs33XuwEjn/tmGRQzmjmvn3vC+RirsT8H9xwf8RSTFf94WitgzzwKpdzP/U
6B/SPCeDpGRi769hD4DUYEFhX1ZUFo+2/+D9hoNNCtw5co/MnSWLxYZM3qXHGMWF
TORc/ZJQseUH0K0p0AYtSSBA5c2OhF0RmVk8Yi7YxDmMmm3ZuCXnZo4HJVMJPsET
fwQJsvCQBTKz6xwQNKh7dMrOfpvR9iaaEoPxmTIxHrBQLFatCL7n8TDpI8Xg3fh+
qhShwGkjfyAfErzz0Z7M0SjKaCCQTCz6A19JAVg/X6N1QBeq5iUXMAhh+uW64W2l
jKaElpPVMcjhdRqyf0uepya3+g/fftMRl/twgxNYDheZ6Ri7k1JzmHH1r/Yj+E4E
sfErIA21uadQZXIb/7wazFPn2PXH8FCw5b2LGf0LP08/TB0BFFF9PxBXWt+9xA7I
LSqvDKvKPwnzwOP26VLgpeH8JyFb0Lsws4m0Db515HrRnUuVWvkdL4WljWVBO/b1
3ChxXRme7taHxx90rR6S2CYB8Dl4pQco/UmEPEiltMydBYZrSAwHA/79H4eX0e/U
rbCrm4rtOKSzXUSqwXU1QkyILT5+l/m2WIng1duOv+oHxM51B7LQmjTQeuUiuD0a
gZ/FohaSBqofVOa9FoDUkWOob/c0YCTzukdjN2yiMit5ktB+3vjPg/zv5bMFeM8V
tv3pG86UhJ0uC6B9KrB1U26CtguShwTEDRrMMCMwSz3Z6qO25wFLsDV4StuWr1Dj
wtJoZehHkZ3aSRlrWsihIbCCJfdXMvG1oD6c++0wmQVcccjdr5BOanAqKU1LA6Mg
Cb4Gbx+8b/J4WV9hxZ/XhSEEWTmgM0bP5Nyh7AEUwqnBX6irkWt7jR3h29cWnEgM
rn7JaYaTYYf7sQYn01zBE/1fNxsLKQbV2VADfhgi0pVoLWFBp+xiceJLe06b/cL/
ipqtvo/ZVJwh2qDnOGTjeEkyB8azr3eIsRD2VTw/owa4xfTlHl1GYGaJgi8aHEQv
UMmghV4FSjqBQ1N8IEOKVQ47iS0ewCbyCyXLprdeG1Ffrys/4V9wjo5bDPN3Tc0H
KWEmja7Ynh7zeLdRDS1y0FRiM2J14OO2scBrdasbaSHuePp15XnTl5Lsldh+ycFw
FxjyJjKZ1Mp19K3o401WaQNolj8lye1PrNd8vFSF0+XvLXt2NxcwWawiyz6G1RWq
QGhTEksu8OpDyHgZELmqNYTJnmnfKct6buAS37/mKH65mqNa+syoahZgJv+7nupD
gFrhJyEH+5BS7JJc67L8KzGdtA7SSEnXQVxg59EJs5maEZKvSYb/ibnxXorZMm+L
hQlTleMn/Xb3Awwy9ea4ZegAnyLh5m6oQC3Y4dDLcla6vy2eLK/M2T1B/dnAG+zd
tefH8ziDX9Q1eyat8RFu638igyaIlJtaK6cXxquMisPcBOAd+ZIfUFuBACp3gIlW
cVyOo0ii3F5KAxHnaH86MmOi90afwVaBxEOoeDR4Jcpx/YzaxvcnMwEw/JjrJjMp
PnFI+ihldpMMgnZWPPEqIqav6hTcFBQ0aKDpTsGWLu7Hz9zl1itvp092dj3OaNNE
kPAytwhHngy8ViEkq/Hz5DrXsSHr4NBiDj1/+C8yRbmVyc5/cctT2CDpp6hWxta/
8Oenl3Jkf5Cx3s8mhwsUzkgkobbANmgJNz83bQGa8sxTak3IEniMcQJ9jH6UmwkD
iGDu2gGq11LO1fGZgX4d+QArvQrj/g2gy/yqT4pFZjFAWvJe/Wh/WcD3pm6Vt6eB
36aq4RYEWY32s53trJc/YY5d5/P6A63VVQZgi/l9WmJKSFJ22OEJCWMaBTT8HVDg
VlcA1awbOWWTzUGnXGVtZj1FCxNzBES7PTvuY2RwLCRPVcduIMCzvChQVVXiX/AM
CTDluwy2EoW0FNoULE/4j2mebS+6+uW2InjrlkGI0hLm32cHWxUcekrmazEqG9rG
u6oCrgbOiHd7zKJTDKl4o0uIWEoTI2yTaJfanZVs+YGxMd/IeChaZTnfNu1PjvZj
8Yg/73eD4jucIzX0LptxLl3JALMqgKC7RhVoKS0//IGCdE7ZUroHJfUuIj3YQolI
lPvQXeHzimedEFy0+mYV2dC2yuwqI1gvkT6o271muBsqScNCMxWq6NiZ3cC9oQDX
6eIGCbqW/SFWNF5o5vt0yE6wPm0zg8qrSyEr9oiwmKsD/XvcGSSR4Q+4j7Q+PUkG
9TWfcUGM42fSAt8JOZL1gm7kdilfn4JQXiGcyye4GxT0aFUOCqJ3A9J5pzE3jWEI
Ci2EP8XaNA6xoTmHRirllqo/Tgq6/WxVgqYu8VLhfC/4BdSEhlAa2KTp3K9SIpwB
dBsa5QA6YN2sUZpp7ehbdrrlHoBmCNXyQQrvn7HdL2Hs55AqcdjtznLZ7yg4n9dQ
Ek3CHoX/ecBDd+bDNXvs4o/iJuitspPhawc7ANSyKsKuZTwlfvOKBf3FFw9YsTyn
9HILk4CcuzGHh6XqPS1C3/bTTuEQe67t97HPs56Qxg0GIWh21sbSCWdfuwTpL5Jh
fhcbKOc88e8WXx8w46tezlli6FHkdgDHwEp5Qyu1XQ+Qh8FO3I5QdZmzHf0Q/vU2
y1itZXuu0yjI9vtzGQbSmWVR3vObGyIL7Cza2r/MgJVG/VCa7L+wVYkg4xS5tePE
iskbRSQdvk1X1xQ2IQlbYuddymtS4gACv4b4bI8zvA4GN/fY42z33KIj/1ecZ3JF
0GMa8xFpkyxA0HPQXoViNLrAGPFIiT8DnBinCTtQULAPcFN4Hy9NghrS8rMx5fuB
9ztkE3arG8DUaX4nLTRspHk4T/dR/iQ0m1v7mgcdQmPBHgdOxEqQEo2gG3TOgrxZ
6Fa5I4kklvXm0NtYXTcQIvMIacr5Vh4xovSLeV6VlbJrfqBKQJEuqzkg6AYlUaHk
6qZ3IDYpb1gOd22Av4p+rdRf4D1Wnilh1xY8rdy13Jg=
`protect end_protected
