`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "W-2024.09-SP1 -- Dec 03, 2024"
`protect key_keyowner = "Xilinx"
`protect key_keyname = "xilinxt_2023_11"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
Swtk8rO9qR9UPhPGV58BalPq18w6eUfJu4ZGnbCJ0EO9Y1unhvoNFBjvzs6r1cRa
0tLMvZTkxD+OvOADNvbX/NrUCsVcJfQMrnmDbKHdpYyXoGYoYtUEyAIXuUXiXycd
bpzhVXzB70bvGnbH6SR8IZvytyE/csIQDSG1YHYlzdxAVxrEFmYP3RqVT2eZTwvB
L6XZdjuEzY9bDfjMLdzivZDA59pI3wMWmrMzhH56sJ7pzX7Ox/MjR4Ws9KKMXcbr
cZ2YSsSE00UHxWktufaDq+Y/v359DqPFgUcB0y+vpEkPEeF+kZmP/x0DudUlkUFJ
UZMERI4Q8X0oNXzm1QZn0A==
`protect key_keyowner = "Siemens"
`protect key_keyname = "SIEMENS-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
LLOlybPtxyKixOE+8NYoTnyqcqzohGMn4B42R8Te78ploRDF7X3eg9uQ0lbCrQsa
E7VtBF1QSbkC23SzQLfBfe+unUsRZo/Ww0J9XQUlrfoygKWD5c0VO6CkMBS8nKlJ
4YWWGjFUAKTvs5kMg2s+LknUPVb8+qvsamquH+k0Co/IiUsBYboX6wieDXRzadkD
7aBAdyKK2tqvpgy74WGv532ZugLDASTloRrX8XZCxu/Pd3jBZcTOupcSAoP8y43J
XNqx0cp1uTuqZKONSwfBbYr0fcX2SZvtcDok+B6uOFtJYjtODiXk4ZXoIx2tC80l
bNvtW0yl6WvMsoGIeTpZnQ==
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
E7elkMJnQ5YQYUEFRUiClMKMF98+tI9TfUsebkDl4aKCXVLRpfy4KM8SJS5QBalo
NunqqDdE6rc/4Pi45BKXfk0U64A/0SBacO7OsNkkeCtU3TB+iWSCuUHHp7hGN42R
bAzZLznHOceRohIXheSZaE9BDbyRgbMrB6Xpebng5Yk=
`protect data_method = "aes256-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 4928)
`protect data_block
smhRAd4NkwZC+3Gh3VwvgqjMpw5nssYQaX5fC/NkjiULLmyXb7cXOr7QvjOyqZLY
gyb5Liy+EeHxQi0V4BaJBLQ/F7ovLqNYjtIkiXVKmnM3Om97oAApi8ABL/l3qZdJ
1UqSsYx962i6CEP0k1z3jWyIq5UYb+ADy7OFrtIVHM7vICKoBnXvIFPjxf+20IRX
4IulwHLhhMYX5+wMvzPYb5NZ2xhhL6uJ5IV5OiR1vSx7MAD9LmOWHuvDtSMXiIRK
2LSdIUyi+EVG089HgA4RvkupGqa0N3c5Ix0CWznCQBn8s/NHz3dTjXk/PM0nI3mz
oGIa2b0LzkRau5hm+sGPthRkYAW0rofP0vOJs+CfdRe2dMALe0HeINexHKwu+NG2
3o8m74d27ADYJMsxh+I7hdC1Qiit83YaLv8qugfhqHvGMbhfyBpebVZgHmRjQHsi
U3xRV2t22nUqRHulc914xF/lEvoJ8PSGaqsgVcClUQ0kw7FwTT0fqBy/aUoKs7ZJ
GPYr2+wfNuRyFSLer1gxE5lmvU6AGZHQloDTSNZwyuTtqr/rNCiWC2ZUspHmfxJS
rU43cFw+Tla/Oajq3snO5rKxCCBFQFHMvk4UPtG2UcgD2brgDsVSyTcafUuGIVq1
6fAr2N+X0U+p8BsFAhgXik1S40nbnXnN7iaFZspsRgh5EycADkX3g4ybwA8Sjohr
AowHQv6H+PoY5YlY1tBZKwahB0G1q1AVRggU1XKyFsWzc5BOqhuzLc7Y2qy8qZ8N
Ljf/lLda5o0AxV5FvcvMSHSgq2AA/5GXfffhzEeOZbaJFPQw3mSyqXVeFeSs2PuX
a4pjOwh5GqMj4F5dlGS7GUPkOxsnSzXjPPzrRgV4OLvzpQgslAk1ic9hiB8/HlWo
kfJlAKYaQPxWiRAq5Cd8ZB5dqWNkJu+npkAnPBQoQGX8/PBihmAN2J8JLNC1/H64
2GM6K0P4li8TWhKZ18plD/vsRwa+vSZVRTA6xhY6MPvvNQEKIQb1Uc3nGvSxkirV
j7hTJXaMFc+36G83a8rVcJ6uxFjf5K3uVy4lHFN/W3Mfsw3fSjo86kL4tVX2fbse
6cY9WLMw0JKPvbpbZc9y7AP1NH0dXTRplCPLuqX3B0bequhRqEn6Y6ug1AIuzGsG
IW3QisHJlAac5v4X2f420PT95elZ+9tV7N6FGvFoCSa08GV7qerwY8Sh/dDjFT8F
J9Z+Jj6ySPPHgTwr/jKUxo3zi5woK2J3AogRjTsxaqd0pNVrgtyZdi3NICjI3z4Y
MIyQ3RBWSQRYauhiKw4hO2t/F2YW97UCb6dm9jAao9ewWpmKxwwls5KwSUZEJxDx
p+xSQuRzcmSEHIC+epGQwIyQWBGgmU1WK0BOjhl/8GvcAvqJMVlJb5/ioobrOyV8
l6k8Pyru+P9QZ1a7gM8FqR6oXbi0VeL3qIU/JP1ek89OZjp/LYf3titwaYRhPNKb
JmOTDODefH0/smS4+kBgnRza49wv28DzfUNLH81KxMjs3h5+yewb15x3RyfoSrmk
a53PbLcymf78VplMFZXpYp82cvJ6ZDz/VfsF2umz0G9x4Ds6M8XebC3zuzIsKu2V
eja3HvwKKlTFuf9711rDQtODJ9VWc6OaWwtw5yjdRRiRKCWp45SfKiOK339XlSBa
opiGR2VNCR+Sp+6UZlF0Lo8FOe42TiDK/ExWuX4OXzDUdgB9ryowR25ZpoXZhGq6
47UZXxDf4JhLHNy8AtUoCOCatGRsCeb1NS8uyZIs/RyiR/kiLZbRsHmJk8uop7qW
CTzeqV2H9FM0JK5+qJow9d2RAfP1U/a0pFTHiSDxlyFq4hxlyPd1DMZuMlMlhrYQ
L+vAXP/tEoDQ+7jGA3v3DwIjuJfxdBMznZ6pBLk2EhfDO8/wo1lOcL6hRKAxcnLi
pyYCRTAJC6ct1MDCaqlsw46KrjdIA+mgOPG7ZP4AsueNNKdk4JJsgqkdWfwfynSw
nPP9mcmh87xFeu1ck/z7tOo9jjVcXr8RB5G86hQVtQyRIb5v1rRVx8pBM+twdkbI
G4rUmPPT1OhTHBlnwCwjCPFcTKjRalMT89F15X4GR+CVGh19B17GU5Ne+CZNdVl4
q+aYP6dKch3eSosVWLlKJpgNHMfUwhEBej3nZDG+3cStRDz4wHnpEBafkGUVda0p
LnGvMqfrYEn6X27lm8aF7JyqELgq1QbtNEuHDKeJykf1ZDf4q9I3ITV/D+VUItZN
R/xpZHjVd//JDUcx7zDTyUVIhXa1CcQfwnw79UQ6uN1iiOxhvrtS3AwzKoHvakap
G+YX7UFNXY/KQcyv9VWaH/eS2StUBX3KvYkTc7wW5OEMC772IpsLv9GkqHsCPMsn
QJBtt8RyF7Iz/5c+m5XTGg6Bt8IJDPZpioTb2RIw9DbG8izwJ6+MbLGUv1XNLDfl
3urzeWexDk9Nz8mBwObPxxJcXSFjmsqZOMHcoTwe3tebaXE8rxW44Lxp0pKWV/B9
JSOJxlybowpKdk24KXIAaMAC0mlS/THcbtvbaFztGti2G0cAxVrTtZBT0g422lHq
kU5/QUv6nUq5efP0uXtuIB8h62qpN2ZJTjnP0Ila3W22iAmbawkx45p2Hv1O9WVF
1bdZ3siFiGXWSCMlhsV9+BQVIApdbFljM7ZXTuvSGdJWdr7BZRs40ZY2YoWTUjut
7y8G4jma6Gsc90tipfT9Y7MT3QgSkf72uUhxPq33JWj5w2JANcFeQcoeRpr3OT0J
wyUihARkj9QCvpAjJnLNyr7nNrEn8aSFLRIqG7Px9W0IiVNOx1sx3TDJq/ayNTtR
817ybuXWCP15S6Ds8U5QMWlIKpqcw2o735SXXrBYW4J8D6r3aA6iU/AubVwJQPdy
vt3wwkT4Fli/La+BdoYvh58+2KEWJWuzfKAH3Aqli/JIis+gK9lUnYgCn/mtkSeQ
SnMlv79kG80s1Z2oWASKeZVFbBdiMp1QQQcuqk9HsD5kvvGYzmfMuzsSilrLWtbA
NOJgFDWsmZB/F8gCVLOKyanYi6a/canFxFy5wlNcWZNUeI0Dxs2FZe0VJgRFeeBs
UyBgmLEICzz8WagbWXBh1hAXNW1Q9G8sl1hrdjOQ/CeYr7eNpiDODEmGt1Nzo90z
ihm+hqyb08/bQiV57M/b9JCpYyIgoYDDjXriFKBzvY/TTOgzUwkohps2gJ2ef2f7
VvO0upyKh9j9QuRaTsG7LcreFZvowlGhetYPB7bLDVaSF+WwLpZtMduu3Gx9cXjG
O9Ru6RUMklB10SD0D31oLui5kBkeOsuxXJBthJmbbuQwToLDCY0+aj9fGz8IKNmL
5b1Vr3C9jTfdl0ygpY+/kET26mVabXQHgf370aoYtMbigjyKmbg4Py+iAW408vIf
RPciRTy8OznmgmyjccdGP7rxzkCN9sJl1t9KOBsnWUdaAlpblNrnRLKS06hv0K8N
EdPZyi2ZRtdMifncXibNOfDvtzN46F2FPNooBUow7a4QKZXesDgfAPbvuF4Dyi2u
SriVgQQjh4oBRSdzC9Ds0bHD3Xc41b8KSdBrvJ6hCvLmj4tg2aWgSgyOaSooKwyx
w9TdQmir9bn8OX/g4nBCyA8srG6k2UWIMPV8MhjooLCKandXmCLuG6vQlzAs/omn
7a43UlcHzQWItnfCF5N7wEiFaLYCXsaiLiBJV7hr7/SnuKUu0PfpmXt5DAEcDY0I
6Me1Y/k6D2KP0uN/hkDi8wMwm3COU4L4G7bNoItsBSME0pIeZRM0qdoDspX0mfYf
g0B0fxpBRfpdXHpWZaTEZDzHkTxcb9d3yVDtAFSPiVHlIvCAOInEeK/Ept4+ut4r
B+jCiKCpXzb5nb3rdAY6mkJIul/QzZ/ARA5zANCJI6h9pjL4uAEI1Drtd248+Idh
OU7pM9jQRhocLJ5aOcn9QQ4W0PTblxhCFlS0rWEMXHayM1woFk8y27VT0v8sqzmV
zq8EDLp4yOLnvvK7P+3CszyhfQyfyp5+K969mM1OB4bz0XQZX9vrUY9UDY5YCyub
xzegEY8N3pJh+8vIlKvDFjAKy0PmDyM4w7g7LVRcQu0o6DQ2HJn187pbt+r3bd7g
uc8vcBR56UnFEq2rD3yZ5ydXmi9M83WvGpTlhkglk0yGeYgE5+r/VCJjsbsF0h6m
0ueG6HJ+29fbtNGJ05OyJAFj92b+aNfBJ62ZRu2twcTmbrTfwHXBjcD30GQVayxk
iEtXOvCTdXPcma/ELhSUiktMfvItNZmT3lNgGvaiqGaZrYSQuOLLhYThYU3aUGhF
VZOWl2TZk2qEw8gHHS0Eq0qOceZzKFJF5b7651n/FqZ1D3jHgwncgjCq3wWF24BP
QKeGP4rASmZRXcW9Tycrcq9WQPBiqDFVOuOKLAbj4L3zZUrVfBm5SnIu+uzN6F7r
JzRsvNTVziJ69fQ3Bf08Ka/0y95Qi673lFZMWRGhXza9SekHMYwgGKia9Ery7tG8
sQMuWFhtFvVuwUGrq76m8tyvMQbO92n5uf/dpee7m67HDWJLXZg7DCRoEZsM+Vo/
yjDus+cqINd/ZHEj7t5K6KCtEDJtkHR+9Jv4jdsU8eXJ0KtxBftdggrSb0XS55EN
JpcIGVwGfqLIEsDSsOmrBEjve3cjFF5QAQ8OXq9+TirATugmwTeHNYEYoB0SUakn
lFHaLR2R6N2UN6paUtRbyt+tLpmR3psr6gss6jIknFHNPiQnnoJJ+3+QQuHgfjYT
U7uu3ocjUhQhYsu8xhWvrF4v6h07h9E9uULwDzH/l2kLyAyDh5zqCgUrxDbgfeR8
1Al95SsEhrCI68xnleKctqVmhmoD+9iBwUuQaHCLliH0fEm0S/bhpSp612BHOjms
/MRvHgr0anQjOQYhD13L4pko34YMsTI8oCNqh2c48QK26vCAerUynxdF+FIRrtoH
NkocofB03KWcc2rV4RKusUpCZ8+KLJ1WDnxMhv43vkSaWdCq6MIvOi/9kaCIhrLr
qRwpKBWZ4HusC8EJR9LDFZO4KlWvGGH5d+t85ozyKmshIvGp/shi4brtZ0tUGCfx
DC7CqtYqPDUOCtfgPIw9X2+XBOctIsq/LPf1pGCYlF/42MGNQvbT8XuPn5DnOi1h
tf//re03fn1LaH9cxWF9dY8k0/Q9MTa04j4Iyv8XJaHkkU4EfPV7W+Fw8PEmXKf0
x2lUJJQ08GjOyalrswV9IEOfsDxczQNeJ/eBd0hUO8yq9K80KY+0FBRVTXzBAWkX
cK7YiI+lUiOImRgWUGyTtBwpivCFMFjYVSzAgqoc3Ewh4jpuWFSB8acrDjyRoO56
8SZUNQIwNH/Um5bTkjZAqYs7jHq/qeYKbL5vMiYvqENen3xl+dPso4IeYgD3Yqfk
TfvE9NG2a5ijzM5J03/uH8E8/bHkkhzyJBrtftnX+YhcA/uXd9AT9TDn3Iqbpy5E
vgyPsY7pLC5J0zT0L114PaRkw1NMa0EvXqP0LefTIE2BOrwlS9mW918xjjfxcGf6
3Lifzk/6+i5RJFuQT2pouK78u6bSmCPDzKaPEWRcjx/XKB7RRb19OPuqkUHVJz9b
u+dQXpEKi8u5lgDVTZBsSBGcFmi7jt8TZpLoOltYGoQbFsarJlpZnAHLhCbfS9BB
h6zhN4F8UQSO0C0SzWxEkEiGHxPeMDMdPLfKxP0hNBhLgRk8grIOqU37aAd6UBPT
OE2XAt/GARUcoPcxMm3Q0yVY7+/IzZ43oSC0pkY9XzRvX1XLsex+B2pgJJESNAOp
8u3gKCSJaJl+3K6jUDWBDAgmPLC/M0jSPHGuX9VeBKIEFpxgmOQnAKsA9ghCxqu1
n43zuKOQ8NLpz6MJAXce/Bbbp84v1hVbmgUf3TI7X3GZKWqOjBLma3LfVDy0nBx9
c3iMzEx6Q+lkfnHjotlMUNGW5cFZkhfLi2oLXzchEEE2UjVCqVGmRpWtgmzhLn+X
n5Xluolou3OiYyBNI4mlRDQOnuxbNVMjDBYGzLt5fBlKIJFhP3AVWjk35mrlTchW
VbXkYciFuBvtcMMDn3XT65nC1p3sbMexqQX4v4yQtuctNYJ8K0SP9Ugr/3aiFH9a
3MpkXLpradCgdHRLMq+4OC5gRKRqyaTTmvrwSRxdwW64DxxGgqv3EGHnqmlfNDzj
3HKBkYladgt6fDhZ7QcGkhQUBzNq0HigKgMEicCBuqq36qNoDN7Il6/5jb1RbaK/
ayKRFzsRv0q3j/YRtjTqwceEa9fOT74yXnYRN0s7nC/TRVhkhWesPU06fq+nkLIL
nXekUdRXU7lY3hPkUDcsqnqr3A8G/y1/64NktDCpgms/ahEH7jf8txw05MEgMLUA
6nTVZ/HJQNOBo/2nSfG63IhJn6uw+Rx5QZr973oK9V49b9imBbb67ottgVZPetXf
MXUEp3/CsupDjzd7OXeaHDP3Sln6P5yNYpruoPkKsplSTSQiUaCXsuPJGpbxhH0h
bvAaQCeUB9pbGlJ2o5A+pfmb1UJC+8snhDk17ERhX9HYFvKSaAVISsqMZ49Ua6DI
OzHiBO4uEufNu1vK1xoK9oRRWoaKSPvaA7PyRXMHxCM=
`protect end_protected
