`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "W-2024.09-SP1 -- Dec 03, 2024"
`protect key_keyowner = "Xilinx"
`protect key_keyname = "xilinxt_2023_11"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
Vi41zhdb9xSlKPsMeUX17C+1I9Fy7EnxHSQUY/YvqIAVAhVTbcK6xLWP2SFy7nXP
O1neZC04stKg02GQ65g4ZpDmVmAYWW389UhggvGRd5qqLRtsrYoknrsCn/D9htRL
qaa/zl0ARkow6p6WHFj5o7STJIYYzO8A3hnQRYkocmqLlhagbGwWHblTh8WdjX46
eBxiHvDt3ptY+RdNqVRRlSC6jmCxg7L8/ltsu7HITRkDCn7dQL0Mptkxwi1Z90Ps
C82pjnJ76EeQ/1Bc0aIojVgI9lbylUq6+9rRPKL8aMS0RHsZK+1UJZloerH755/i
QXpGUtCHbAGfUPXqQmVv9A==
`protect key_keyowner = "Siemens"
`protect key_keyname = "SIEMENS-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
uSFJBz4XOGa04uZInT+37ffl0xGbJfVY7May/+pDJhFaQ8E0j/vd36k0pS5m11c6
jq0hx1v2NmiZdT7UDyBMl/OvJk1GIwybpaA8tGX3IMozWye0DQRpQt+e9LMZcZHP
V9DGTyjrvpA5xdEea7Y9USOJKYogXecXySztsbt8BnM8NO0UpcbBrmc+QxODQqlq
P9iAK2LYtHXLqyoaviZnyKt+QBup7WBjdE5pzRYKrL0nAFbf2RQd/f1KPDHOV8IK
WlzDQqbLz3lThyVPZ5gcNqTQjQh0meALLW8bK6LJDMPMWotr9FCxh49vHuT2a5lU
mWRFk7YMTwr3IyV5rk1MjQ==
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tfkELvHGYNDhRH0orfGTCbswZTVx43UisgKtQIF1Z/kX6E5kTt86kIuO0bDnR7SG
aaFozpNv/BMaPjxwLnkcm8oQW0NTwynAxR65hX+BRkJjvC2RNoXq8tnlIns5R+Os
XvLUJ+Rvfm3qiL3+MacRs45/oqmXbYHOd7GDyahVrZU=
`protect data_method = "aes256-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5024)
`protect data_block
fGZDV+Ab8DFiLD5WvQCf1Fcs+aEoY6SzeEZlATOxubvU10sGwA2yaqUkpK5gTOA2
3boKvKvhjf1aCEC9ih5D3egoLlMhNDXTg4ygdYimJug7THsYN7pknY4K8aO1AD5K
CTIaa1uLofE/eFxJ0/dlcyl7Uz7y+ugdxQlEl9MC10J+bjPy6ilON/CqF/V0g+OK
mmzkR+VbUVT7Ucs/eG+cd/kYSQoDRtHzDpV+5fhJiKBU50KCc38GvCEugN7IBZb5
3AZpaQe6Tfk8/sAW3wK9VWu8zs7VOEjTayJOVI6vErW1TJdvbFois9w1jITWGeQC
KVrHnUm50/AZVdLaeVr0sLHAnC+GWMIFT7M3zA6zjCxkAEWzlwjsbe6tJ+1530wk
tDaC70e+jQPpJC5qvuqQdHaI9gEjTzhx6Iu+ISDTjmRv6xaDc8e6EXMvyqOLd2KG
O5qNERK79LwRV0Bw5r+C0dBZ65XQUpPMXHpHOP06m3cYuOVw9MI0yITfTpWhW1VK
hJrrfVXvLS4aHOPH+Qso9JLuSAZoWzfRQVFBy9HyQO9F0uK2xOnmGzAWBYWnEokm
tBoLCT48We6Lf/PcSovTjLSyhgidSCQWcux9aGPa63iaI/abg0d9VOQF17ScJo9f
DnM7Re+XKxbPbvzjmlIG2fBwXyidVijzylXlB8Rd2RzbKwmgtPqPbbczF8oJ+fJA
A1x8xG+DFbDOtRO21MY1y2j2JTkLT7QkQVl9gaRrhwcNLYz4DvTq2fUndDuBmVew
Ymg4gQYMm27xVKnfJEa5Y1BUIYAI6x+nzRz+NCwN2wN1n7D+pRPyjGJdOb/4EIua
o91YQXgvZEc1K7yFtUD5tOoiaMkmhNa8AAZFJ7Sc8bL9c06fjLERpIzgWZxl2Jdw
SRrpSl06c8pygjy0ehatRxU9S28BGAUTEO4QaI9SpxlqxWR9pPiGJ1cmgWIQ/QRv
2hahABVVbZRuOaDl6+HIlQSu8vktnrLYM00iUk8AY5JAQ3JV8Il90ZBrg+njoGli
mSrbHBKz65tevckgKr1wPA3NOvs+yg6mFj9hnKRtTmDOkNjmepG45Bx9DBw9G4c0
tj/WaBgiGoubtqFsSnc/xyTiUkjvWxcki50GuJypU+aP78pHuYpCohTfVxCKwr5K
OuJ85s/dVleWT0M9p08vI4+LBlzO9bqu1Gd+x9o4VxLBVKI3ajAVfGLJqP+dlygE
AIzmjQoj53jrOUZDW+NXAxvBLLkn0GSCFMkeU1YBa6Aozso989DI9NbF7PEEQjar
eeKytR20LxTKFjrhjPUp2bw8GFWBT87nYvpzEJKe4MpSrQRriid2rdBZN3gcmfiO
jMwUMBeA3aEPZPmN1nSnVOjjtXFnC9TZ29NZMC+Mqr8OPa0KFwwgW9hDWk3U5uXF
JUAF+bpWzbWEIJFrvCzf7yMGj7Ska59bNhJ0kIa7p0oogXlyF055vTuIZKeD6Mnl
h35uZy8nPOFdMIrxLP89ZC/GjfjaZDTsYzwY1VBRMnJz6gMXYI5a5YqshrbMTYar
kDV6TqVMGvFxAMXa+ODo/Lu5LdLS+CBLv3rB/SQIP7Ybr/R2qKzAy6JAh2PmdgIa
u/PBCMejX/FVmy9a/vmv5cpo3eJPhb/HmaiCrEul0dAs9amXFvcN902TkA33bTxI
t7O7Hpeua37dyZruCQ9cfGHv+bkUnYmoglDneLciRqnbftgKZ7jZURsMo5ai0ZjV
Y9lDPPis6HqpcxHFSGT91GyjuvAq1qQFdhC1KW/e5lbixVu2OY9Bwv0cXSEMJEzC
djL5FRObDZ14Ebg/uSSZ6qFQfxHQwToi+Iem37T6fDfaM5vV8zHxtv7wU6GVKKkQ
Awftnw1chkFkZb0bkudK5JoEradujZKps3ZdtFZUZr6ul/crPoPCvQT3R9U8j5bf
SRTnUo+Hz7A1Y8wimZMTU90oQhBc5j/5pIhNoJqh/vy9Qf6xki3heQddMAItl4Pg
Dt3MuKckr9Bdm4PHITD8AJ2scVs84MMxLlQb270XF2MdLTp++Ugw13DUseimSeJx
lna1/coP51BuQSkn5RTJllAGbov/II/8e1zwXzZ34OlxpXUk4+0k3ClmUxOXUBkd
NQie+K0bfrSzF0r794vWE6npCdR4Kyda4zdlQt5jpKVolYLfKIC5wfJUvsMdfSLt
URVWOwxndsFCDU4JQHN+8IV0CXV1NR3Qr+viXBY0ZiR00kgNUhNQZb3k0WFoMbJI
bHlbACuWyr0sdECBwZSmNFNljF54aCXvICVEkWYVy71wFoi6/ztR3Xh75p0OiJfm
DhMpLgDV1qqp/QapdQRr403N+yXpZ4z2cFZo2xxs00SSzkwH5uo1nxsXkL+17CKw
ZJy4QonZpgoP8GOI9rGCDP4u3mY+snNLH1jMpx2Yaa5dxLzbJYHFqTZU40Z/6wXb
7xU0DxwhwiOsV0/sr1eNFh8XktnCCBHgTo0xCe9ja+tknDJ6ATOhN1wSu9+pbS5H
fEwJc6hWJ+cKupJjtUEAQDlF4YPeMxvD7O5M+UMUd3m1PK6PiRzGBbuTlgUKjYJ9
N6vhKo6VwLrXaeXFP9vaCFee5qJKyPBiHNHwPrt8pXGO06Aif6ZP1t4+D92fZWKv
C/m34AYcNxBW7+yK6COA6ksXMe1DSY6y3EuWNz04ePNDPrKCb96y18370WkeIuet
zKUPhcRITgWYd+EmL4AmsHEk0ItERmfCGrY2Spo9QU9BoqWCa4yFSdjbuxXrx2E4
m56CjjTufWKsCsdAYofOsNFo2ZKNwIOMsP4MDVjO7oBbwviL3ZHwz6Q9UU5G7RmU
abcC+1DG1YZLfeI0l8FCJzinbvXb5UAgCjDDwGwdKTr881W0CJkaXXcQZo3A25/w
+uO5oTzWrp916T/hu8tnDycx2lVY3bRYlyJ4M4+W1+YR8tzjYq6BRb47zo5qOrsY
5TgAPcMTfzsN1nC/BIGdBhVKY84NHpOWXUpjCCkfJmch39akEVTQ0QxazpmEAU2b
tD7vn4nBAyRr2qRdeyFPQugjfa3G9C2ukcUgILfrLuxQq3la6oCBByROp4sdLkKz
d2cZHoh33jgEzTpYPYodXz1ncZlCe3SgiaFaBjMff9rTLss1WZP4QJRHulYtk0Uc
4J9DVl2+8OkIik4Gn3iPECAgihOeJMDX0utLwZQ7rV9HJpWEUWlUUegiGDPjT2z8
7wZx3WzH/cpeoGGXQtplx6vM2y/ZC5sCBPq8PC1Q9JgBVWYvlJMdiV1pp9FXTNyP
9sMbHZOGPlSZdUcDQuxxkDyuI8AHhbN5JjqVCiHnJAwaDL7aTs4/bsQNl3GREZG6
XEvg4Qkbma7Na/KM2E7T422oI/9cYESQsQNEwboRUBYIIZUFo0iT3KTZc5erMxzq
/RgA958/UrjqTXPRwTE9Kn2K0IVQrzwZCcK6IydYD7pMGX7GKEvb5RZSBksoAxq/
n2E7lzAw4mIizndKlq2wwyLwurMnlEONpXqcrsCg5EeEn8g2RwhGXyouLJs0MCm1
nyVJ8/esQFSIb2nIAyDoVd6eoUMwvfe1E7XuSpmucez2cMCA9hs3wxLiuX1/KrSc
A2UKWEH+3xkHqZR+q8MIy1yNyJHF2RHJbpZH0UMFosG4A0oRUHiI7MzViKm+i0rC
U8kylznwxGY3Hfzd9bF351IH5UFRRQg/3Qgz6h4jVw/0tIG8G196oZFyLbQm4zqy
ltXaMBgzLPtiEwVT4kItOuwdAZpuN5cZ7pB7W7kRQ+MIGRrHmmEJpeKK1rkvhcr2
uYbkZHMMHwa/Cq5CvLUCIdWGMkZJieoTp4dE1lP/6Hidgg22h+/yomqXquZPga09
sj0CZ7Bp2aTSy8sRJV+HrC+pqI1W3N8ziJ/U5+F1Yj5Yu5wnXdF6rNp++gM/H2Lz
AzNIzSuUYqLLfE1jSGrc+nHtrvkesAY1XUDA15rb0p6RVuWrS8DpjG8Ddr4m+5OX
Yvq44BX3X+3tP8qjNQwTp0PayaR86G8ZA1+RtOnX6pjAogCIl4k/j0bFOUF4ZhQS
9eQtgKYPxEm0ocFgxM2SCRbwChBebx+eOZwAwFM5jus1twAJU1WW6Y5HWHHLQUXv
/OactWFqoPnelaFyH1jt77TkCqx2/Bh1MN0g6gtCMA1V+n8Si5HRFd2QnJRrQ3yf
9vq+WQsFuz0qZxidAQkg+m9jkqdV6ivdoapMDXcZ8eybUde0exrjqVDoWQX0WQ0Z
XBOyDlpJmbW+nOCz1khVlCcscf4gEakFGh8Ou66Vq+lEd6zwlEj+g5S8daqXm0o1
bvHAdKS1ubL8cqoYOaST44i/Icd1x35afLLSPdcZuxFALs6SoXxot29VK8DYe39P
MoUBm1OmGD8QKKV891JTyZaxfnJcyyeZARqMDj7bh/zmZZxnJBHTcgI5HW39Higm
n1cO9WHT3PvnNNvU1ER517DuDjQYoXumxIVGKNA+Fk6TJ5VqNXtpSHVAOrNSbwo2
rXkYX++Y3zx9bkolko50ecYP6Egj7gORjHbTL2yuoN5btgZamX4qHtUSHetUoDaN
UNgQlVVEZK5xAN0Cf5dVUUWZ/DSLP/WzDIMRWe+edcjISk70kWohs/8UOy97xSFA
r7JNEM1qCisi/x0sWqn13zvUcjWzjR13fqGdg8Ic619Nzg85tqMjDrmOb9rjf1fm
Vn5SudIebaywx2WYQs//JduI6XxEE8ujdt1EX40nQMp8/DMRMtorKpxmUOrfU++r
YcpR826BQyvgkmmaAwhMu6p4g8scAk0uPLBMmetC6C7Hzgrkx0N0yPIcxgis08F0
nEZcwDBH+fTP9CEZOFHne6sdsmIOo2gQ9j/zPwjUAGsWGzNPmANF2Aa+YckboWS7
IAWQg6V5/BZSzPhgx4UqpRjDpWSz6ASrK2OZXojsK8XFHNoFWG81NgPKqb1Ujd+q
QYZBSJatl2MbX3F9CB8APzOKe/6Y+DngsIUcZF4F2f+vc0sk2jmftZgM4Gw2OAM5
YgSv4GAN8ItTg+9x909tVcss6jJvJUZxUitcHZBlYCDTS8jFaFPouUjAAw/Ff+2S
HDqRoARl6ywC/fZ+eS21IJ00icRSZ+qWDUNDVAuB/qyqnWDIWV2UW3HYBpS1n4XA
YSMkjL+43oJA0fnCFXx7SL2fU0GDXQ3XJRr9RuOXinYMpX9iwHaFYxnv4D+HiQVD
WKrDTVOp938pHsQrpTQY3ixvYcxSFAZHpV5ZJUSlKtf5nGXwuljjtYglfulMcItz
pMUV9fb9XGpuh2IeMrHk4ZYdmKy61fPsKFMH7Bb0izO7DQUGEnjCgdXvdOxR4tc1
GP/JdntV3bxfASKrc0paJDgjUrbD87N69VG588yLH08Y6P9DZE6Guts7ykenNQFl
8HkQ28woVtiXOEZCMRQm7KE7HO9Hu3FIrEqSZvGnQXiD2SHDv1ckTy/WyhUlmusA
ltLZEB3W1Jz/bwL1M+DVhaWSRg6m0kFvXc5Lt6DWZ4siqsK4sA7vpiOG3tK57drY
SnCIlC5sYdY5TUbA0tPh/tHRUqxu/r9cXXP3KKjfVfviTYanbgBHIQnC3XxFLyb1
D1BIILfYe5P7b9M+AQVhJNshuhsor13vSHMBm3znPuZF52uwzdwHZMwZ5Ka4vBFG
uaWczHGcof34JLQ/D+SGFK92lbDQrBuSQBF12tuo1txiwZWsuozWkhSCp8FrPkn7
4TJusMlc12KJu6/cBfs2pHz8sro06hEmqc5JZUUNOmy9tUCtl/R2j9JWbAtqYkNy
cVAfUD2z2JDsFkJNldh5liHjKEiEMVnCOP4anJVRBbWIELNXu+MJiJj3iHuAVHx2
K+remrd/RPaog9MqURyCZZEqBqY1pqfd1WmZcd4vDv0t2QkCHwOxFIK9ZXivzFw4
cCA0W/H4fEJ+/JtvqgbuBIHUYCWsE4JgtVvTfyzP5hdHIBFA7abqfoGGW9wg9lS6
FLBQWlt71cM+XDifNXIpEbwugRGizlBVU0TuW57aIJgVekljEg+DOtcAo3VG3JaC
QP4XRJG1izvZge66SqHZrhTfMCA+zvSzqL9NE91B+PJq30gpLUhyWd/AnyKZH96z
wws5/Fw8S/jsNC7qTzrujHkE9eeft36QAuJ33oFX0QNmISoyX8j/FFsOdxjbSjMT
UxHRmRJIizJiCx8Cbkt2NDUUJajVJvTEVjiEEHehUtA8wCc5iIUCrOwYpCmgHkE+
+Cu+MVzOWgzP6WfABKrB1gWwYGWDiIY0PsCRTZalsMlMi6AeEdImAadfXC0ac7kN
aNK2fnvGU1zTe2UQsjAGvQc8arlrpCTmSLAamIIUFDiVPxt2micP2AHPIYH3Ww+0
X1fR7mEI6c2+dzhzgLnMvaGHlJ+nvYQrOgOV0mLG55AAfUBbHobCXUgeBne7oj3M
BrjuYhWdgm5/MPt83KpMX1Z+IYjINGUWV3KYIgXCQ9KTcZ4mmL/PqK9+4lx7WsPb
8bkbuVKXj931N7QYAwZPzYzCY/HA3mRn0WL26fBzfP7VjcFZkxvUm6mMUuXfYA3K
U6oMPFcdlXCqGOfdy+0YWCv8I2Me9Mg5GOpR8n7fK3BypGalx7ZoqgZ36y1Uu5Uo
6uCKsBtQK1pxc6R5vMpnkrwbmvCTJLr1Y08+UZ9hh7TFX1cVcp9gTnzdoe/cUVUf
Oky/8pg0Csg9/6KlNpz/MAexe3N4OnLLkaf0FguLMe8=
`protect end_protected
