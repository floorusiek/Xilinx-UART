
`ifdef TASK_1
    localparam TASK_NUMBER = 1;
    localparam DATA_WIDTH_IN = TASK_1_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_1_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_1_MAX_SAMPLES_IN;
`elsif TASK_2
    localparam TASK_NUMBER = 2;
    localparam DATA_WIDTH_IN = TASK_2_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_2_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_2_MAX_SAMPLES_IN;
`elsif TASK_3
    localparam TASK_NUMBER = 3;
    localparam DATA_WIDTH_IN = TASK_3_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_3_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_3_MAX_SAMPLES_IN;
`elsif TASK_4
    localparam TASK_NUMBER = 4;
    localparam DATA_WIDTH_IN = TASK_4_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_4_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_4_MAX_SAMPLES_IN;
`elsif TASK_5
    localparam TASK_NUMBER = 5;
    localparam DATA_WIDTH_IN = TASK_5_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_5_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_5_MAX_SAMPLES_IN;
`elsif TASK_6
    localparam TASK_NUMBER = 6;
    localparam DATA_WIDTH_IN = TASK_6_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_6_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_6_MAX_SAMPLES_IN;
`elsif TASK_7
    localparam TASK_NUMBER = 7;
    localparam DATA_WIDTH_IN = TASK_7_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_7_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_7_MAX_SAMPLES_IN;
`elsif TASK_8
    localparam TASK_NUMBER = 8;
    localparam DATA_WIDTH_IN = TASK_8_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_8_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_8_MAX_SAMPLES_IN;
`elsif TASK_9
    localparam TASK_NUMBER = 9;
    localparam DATA_WIDTH_IN = TASK_9_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_9_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_9_MAX_SAMPLES_IN;
`elsif TASK_10
    localparam TASK_NUMBER = 10;
    localparam DATA_WIDTH_IN = TASK_10_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_10_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_10_MAX_SAMPLES_IN;
`elsif TASK_11
    localparam TASK_NUMBER = 11;
    localparam DATA_WIDTH_IN = TASK_11_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_11_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_11_MAX_SAMPLES_IN;
`elsif TASK_12
    localparam TASK_NUMBER = 12;
    localparam DATA_WIDTH_IN = TASK_12_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_12_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_12_MAX_SAMPLES_IN;
`elsif TASK_13
    localparam TASK_NUMBER = 13;
    localparam DATA_WIDTH_IN = TASK_13_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_13_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_13_MAX_SAMPLES_IN;
`elsif TASK_14
    localparam TASK_NUMBER = 14;
    localparam DATA_WIDTH_IN = TASK_14_DATA_WIDTH_IN;
    localparam DATA_WIDTH_OUT = TASK_14_DATA_WIDTH_OUT;
    localparam MAX_SAMPLES_IN = TASK_14_MAX_SAMPLES_IN;
`endif
