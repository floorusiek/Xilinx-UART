`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "W-2024.09-SP1 -- Dec 03, 2024"
`protect key_keyowner = "Xilinx"
`protect key_keyname = "xilinxt_2023_11"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
qjEfKI92e6xIYpdrhrCDT6FwO+nwKxKXCxpEy3yA17OZ2WzkATcZFncLh/xbiyvV
WRor5n/U3h3GGL63hRVjaQ1Fp07hHHSXQ2s895KPOgLO8aRgN9QRwdoI4FpXM61c
j2NzAH90+3UGsovMk8yO0bAO/G9T7QlgrHt3bIPptGVl3//JPD9WGeBDqnhLnbZ8
f34r7itR/h7ckPGTu/OzPSXUAbBYECUuHs8Bbf9DPbav73/KZsDgNDFAPw4f2sZD
S9/Lji8SFHqJWvnbvr/QMRBe6w6HVPXZOTGasUdHoa3W3HXdYyqZOBcrP6sz4dbu
FmEPN6xtNyOrLrhgChzm3g==
`protect key_keyowner = "Siemens"
`protect key_keyname = "SIEMENS-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 256)
`protect key_block
y3AHU1nIbthbxljYv5/yqjB9V7Mlo83l+DdzHvwf8Ir7xCH5XfJgwat6Mfi4Oj+0
H0BSZR5zBAYO35Pl1CwMDkmSDGlnlFl1QmraK5FXgvnyII7xWvXk+hu+SmRWiQu+
ThMQkiFRFCJFGqc9kAPpLDFh7mQVcLtxXCspqJwp3fyvw4rtOM21ip0vnSHUtn5a
yKQ3iPjbQ2nN7msfLNRDkcapFFQXWn9Bch7FPtvSNY2maGL5elWS8/RO/4v14FZq
o5wumlqiUanuXaqWJ/Wgc+aATofRhFBAhAsqU/9ZbAY+DDZFzmXseu19PJnv4OUW
Gu65t+wgjFxxFdIHOPgzTQ==
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
b9pbTPq3xSyfFFZKpRAedtjvYLZE10QYRi2WPlfAPWHYUX9o5LjrzXyguZZ7zoNL
pJSqi4sLjd8+6Db25XIQgeytd7MW/Q03WtTGHWeRLQ6BXCJ0oKj3uqHhU3bm1afv
wDdXHzy/xC5CHoXusIqVe2mqffJEvR+4gY5uKrq2Q84=
`protect data_method = "aes256-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13904)
`protect data_block
dViuALsHLEzsJuaJP+rtPyR/fnpOhqaaARXCTSqCSphMVBqJJLxMXcncVjhg1N3R
KrMwpY6c+XVzxRAmjhzsvl2XxBSN21S9hOLg929ZP74dDjqv2v4J+sZz4LsmWHs8
pQEoy4y6voRGLUPWOs1gOGPzY4PBfG/xBQtMNs6gEKK3V9S98N0s0qDpf5CM0qUG
1pucjhbwgO+M5/0ySDHwLzk1Xcocc4DKmne0lajFt9oIQ6g57B8HHRVdmvIBO8xT
zr5Ox8x0oOmF2ab6me3srmVvunOjupK3clkVLC0zOIjPd1SjbnKcmnZvEARj9HvR
PLpbZtISwYQjr+83CWtywYfrAdcX5D23qHvW1xkoTUhiLS2tkQ1AF2hK7afcaidQ
R9OtH/Q65hupRLLaWD7iauaNWGiHptX+9eQe2dCEfBvDQj5eWSQIvj3+nX1Q/Bp3
RMbJkpC5lS7DAZuN/6CmX/XSlTdRFp95fVbiA7GsMo5Ln7xvEikcYZQRnaQyzHFP
PAgBowTU5xciT9UB9JZix6kkHaBi+Ahp8G50Q7mfze3UsUxDdOuVSt7X7kZDCiQO
srIt6rnWX9+J38e3mes7h5WM5REjYymjrpczcLPMZNL/0Yns5NxiICbKBaieHIql
w9sEiACFspt2/NydDFMYRDaPLeL9KOtgbc3hfizfnWxSYTVcZg8DyjCf1QJWd7RT
ybg9z/2plv/r3Fu7cerS/xll9PPCLBIk5AF0ukBMY60hYaQCH1cuRZvwQzSD52hS
iJzIQgEx6Sku58TKeJemAQOfLCLDEMopAW1ZNzyeVL+ENHgR5HwtA5Z2p/ZDn/X/
6pCEKgwymrg8gaM3wxu2nERViThikHEtN0p1vnrav38mKfzN4dq+gTo8wIMcLSnf
9GViF7qtOy1wv1e//A/9pKH4g2DwZIAT/+8A51ULONysKb/h7oKb+U3s4UBrhumQ
dR3jwyhUCOPyNr+0+6GbTcoD0NWVVEx9of/W6D+/KUPonoYTEqWZjyAFqAC4bHOy
722uYgW7SS1ZZ5LrV0mr2go3uamUecz3VBd7NJp/REA8racJChXHC5CX1SdJqIPW
gNzuBelBVKSh7c0/fcv7OcJvFvikrhxjfdQOyvZE+qPTUW1a+UKWFTu+lWy+isfL
ieNaSqsZwMKu+0xGjV75ucKubncgOcjFNw2FxYlOeQKaNax1Sbonv4DHgNemyFfw
hRFM+Wt81IrqDx99j5r8BUmgf5ucjyG73JT8jemcx0N4WvOGSl1MI1x+giHWHMli
fRmF+b6LJaA9z+V9ZugCyhcJYNKIrQTo3VYtmPhgeUyQ9y16poZ4/B3QZTpkAS7A
anXp5HkdF+eKmsrgmJrOcVtEP2GpyVDPIbrm6XDs5XBF/sWAgmp5xzB2zI2KYENq
CuxaYZQOhO8o3X9sLPNtj8krfVnDMLFSYjCNmBuN0+Rx1D89vDCYOLefmh6GoyUR
XomIU7mHwMDPsE1iFtvNl6/jc6XN0GRbBqsCOZOC2fXxDW8UuyT1A+FDpocURxWV
m1b1nLeRNTs6gKd9SwkNygVJpIDl+L4tVzqaSJcPNxmbeoECjr0PJyMJT4r8l1Zc
Gjd0xBQDB9lTY7ZLi6zQ3d3VtyXQCZ0Z67T6JJKF87RVyUW7aSb3AzMHIwoFkK6o
sbgLYHwXrjdeCAeLgNldpMWvIJxEHitSVhx0+aFhdXQRZ4ngMHxspcJQOJIf6RP0
zNZXkBLI0yFSUuI0qrfZDd0lj+8Ft1whna3w0JEOCKcFbzSei8Twau4vh7VCCnoh
XvR63+eNGIe2zUSNvPB37M4ri/qm4jatVOJVL+7IyM0nfOA1Cwc7DRzb2qcGndWF
ejof1TOvf+ISb4deOi9VarSvsi9oXgwR0N0m4V/hbeD6/dJ3yOi1w11E40yxpcpB
EWirT2tpHIMBnElF9sHw6EkzC1WpRKRJLpG5NLsU2EPA358Z5ATxbd+O3UzOoOZz
EvcIjVnnrupgGRlpWkQToEsqZcZ3JVmT6IikE+cjB9p3Oe6/rC+yPbC6GbaZUXzn
2AqRLnj5PMCqc4DKB639h9M5G5lsqCGRKb7nRpM6IQyJR7CSjojqU1HvmjwE0EAw
jaiDAvjubgQn2hSkboTGwBmwdevisZOW+xOiQBf+AE40Y2HSLwBtTODMhDgoBQeC
X+flgnKzMsLmJ/OpCkUk94vRZT3FmHLeL/Y6RH1MKM+xf2MJpdP9pTKZHyR3tSZU
C0091aqqsnHeR/6UG2cYt3oE5RHfd6nA0eMMKvDHNkjdQc3hNXyzrK8f2tdoRB5H
a0qjPNz7llR16I1eURUb7QSMaaLfEHzW3mLTXYe5g1fwxdOlG7M9Z+2WIaEAc8ZM
TOj4UEHfcKN37y+JMM9P+zIGpNjBLAZOG9DwG20n9Y+m4XwEtk0ekYfOxDjlf8QY
Rw9H7Ls5zHavQ6Rk4zyh1XWUt5uQ/z+x8C4qLPifG2LXi2hIbH0W5Qy/eCg/cpeW
5P5gxQsf2o+mlfsxlcpgdP8aT25564PihcoygVBNXECMUxJPmGqD0FHWt8UnXLWa
t2SlupyXhN2ha69XqflwgN58+JQdFMtld4TuNiQZLLtFj/jeBv4RWg7yE/EWXjS2
h0Of1pkDHunlNdP7NDvgHFx7a49HKbGXZe2aP+Fh3JCVxGk9eH9Td9RxF7LIDu9c
dUEAubHG4/tPyOPw5FqT9POLEgMvoCdFDjIbmsIwvWL2uT70jcNSr6NA/Uxyn9jf
WlW9jW+GDEiBmz8vqLILPFQ0caamZSZMSQuLLVxqE9jn5cV4h2MQid1SE4jFHJ7l
/AFsBJa0klR2RiG3ZVy1amCrOVBoSyhQQZATXyEvXDEOcMeZse78ibIirIyERlq1
MrquZhy8rpcFoHZDc0nHCjsG8xgMdaEt5gwUIZkeaXqoVCNp+4Mv0OWtxU3JDoRi
so7bNHYZ08keDYTbjT8FZNrjJFzH4S2xtqDK38PRqRH7Mf3sXKO14gAYhesdb0xO
BH5mjZsMw8JMN7GrgXPEK78vdkO/cs2Z84pIw7ocfK3lnAzk0rHcweHktFVHiHYb
4VlDaLTNXewb4h0BrE6hhq5B/lQlsAa7Q8V0NQf0uYiF7wszDFIaPvPWtCKMgc57
naA+ljTWJ8j6FnMzIOs7Si8WWNN5kUkRMqvg1DbHOuN7Im1xzdf8I5D2SD19Avum
fXu6IrbyKoNn83YiA4A23QsCqTynPKqvdo54pc17rfUamFXHnCtidCQm6YXTL+K3
akigWOi18iW4xuOWVyCbsBdcyybvKsTzHlwyFYZRcEJb4C8OND/rzXLRvtJbVddG
Ppn+wC7NGTDqIUwZDOTb02jAYE7XEpJ4RuQwW8OnBgCEDa4xuADgqXNw25zYnacK
J6zdImFrvmuFKhjoik37OG5sp5P2Aq5PC1F6m1GSYF45fgYyt53iyFpvmdaun7wG
xsYADQYQraqUusazz3qJlBj9cabRRs/92S7FWO0+dwtrK4s3Nh8PNtdUtFL6VVZk
qPYMc90/bY3qCnHJ/SG4EZ6rrLQIdp1T0q13hxwlLUrlqmJxUids5gouRxA9r/K/
8o9R3pu/F3X5GxGTSJr52YHoc5kuJsTx221wI1/u6/oxVfVM4JPe7MXE52xt5eWU
5lDLC75cVnTyYiUp/NtqP6VOeNVKtOUff37Mbjki29l8aAucRh6m+1sr1tx7Le2F
p514PntWZKxxjh64Wf747lUAY+BAXCS3F/GxQKFN0WPn1M9GXiq2Smy8u11m6cbk
Di0PL7wE+Ci+mA2RuF50YQ8a1p96FeQO0gCIKQ7LvCGe5lFCB6+aKIBA8QD3UhVU
91cH4UoRaTXiXzDaM/qicd8SNy/V7XShjT64sGJfmNtEu2xOkbM5y2mYGSlVhat6
AHJ8vU+13yO4c0dCBpYeE8NcK1Gv8Oo8jMkIHE1PC1UgeKdOIyr3E3jle7r4ZtxY
DmZv0EbKjgFx1LoyWSUkc2u96p7D8M6+CfsPPHcova8HkTDX9J6tXretQysu40b6
C6JrcJaCBujgyf4ikQN8ubk1bMfNOqNwtdXkbE568jwumKNp1QIqOtByKK5MFJwV
y5Lr0R27aOQr9h9Lznjz3Us3Xq2r2Uk1sYX8KaGxbvrFdO34wsN76PE3Gz/1q36g
QnLKYT47NuSGOcn/hnKszgbjCrRoRgLrTWkMqwW8LS9X6UaqfA35LFgTtzDQSdg9
4CW5/Ip/GrysBIMbUz47ZZm6sFu0HL79hqDidt3kXZOvBkx6+Tx2NR4i/fw1P1MA
+kwK/6DPzmY2zVYRXO71yfQ06ZqEIwE3gBzbgOCk1RMij3aNxWe+3IHNHamrhu09
+UYEMcuVN9jlQgERE7K0X9UrxPHUQlWuPh18N7/k8V1yOenQEUxlfBXHsof4u4c1
A7EuJFaZRCQpGM/iGn4MRBW/eSeJs+0kcDedbZ5HM0vWFcqXOmEDj3YI4j5ACma/
4Yx3lL+00VY+xCM2z0ogvbkv87TN/eccbTVA2bv693MpUnCIZ8Km59kCw4gL9uvf
srecLabirWr26WzG2gYFviUDNrBmyBeSk4Efrz2H4FYW0433CtyF6s9wWnDbxtBV
fO6fREfH4XBK8IYbMj2E9dKwWfd7w3sUdrjyU4Hb3VM/9GyOFeEej5aRTzAXVwPI
krriUrvKx61t7v7eg6fcvdmzXKyEDuWrwsmNH4E1g3IqCrLmMPYsgt7XjGDwxN9u
tLw1DXGYgSIeBO1Ea84GzKbUKJ56VWw+ywdPbRLvwEbOVatJofIkii4gcSQwDKqL
4JIsMylUEa7Ov7uNu0Cy0seS60x3PPG1FcMdKe0beehea2Rta1aJ6mjAdJSLnCeZ
CZSlXLSgEKIOf2MQWEB0DSDsILxow02HZehZy1JYeKS+H7523G8G/z3fzJqj2AaJ
kGBmCoKyd8GitZjNYMnpqOZ3IQhn7wybnj5NSgd3HigAF7TjXRhii5bry1svTIzf
wH3N28gen8m5riOXGKupiQ3LMqyPrV0xPcyJoJUIDRJAC8xfWqee4BxBO3VzQddG
bfkzrBhWeSqN5z6UJfP05WMfENpZFDvekcnyRgWru9gzHCvQ5d0MDtzDHcvnaSkY
wZSnwV09ruuaKXxqjBrcA9YaTApc7oRNoATuN7lFY1p+wak4zDfG0flO5ziRittb
2fbQqKuNlKInjlyHEfcr3tRH+yLYr49ylxgOmvAjOEH+VzczcImTJ82+YnAGAA+W
A3weqv0NF3wraRr2bzRj/tawaPQ/wNTiqvnhE1O1dFzf83KZyA5iqdtP6PDOlOe/
5c8aO2x5z8Z/iuLvXMahb+iu2m2BG06fY4hCZuMvGpeS5g2VXAKHUDDF5iecdAcy
s3P/AbGhZ1dcAk6IuCS5n5KKZau96LoHxg3ZK47fNHfm4+qxietJE1LCF4snofpE
6GjFsRXyPtGI8vA/ZAVsmsMV2Ag1oswV1G0Lxy+AKMoATE/gkibucNhovGA6FR5A
eJ98lv8tXlKfZZcEqAAQHyx3bO3mDhjRIro56kdrwirYGhFn0vnDi5cAk81yviar
5NKYjOreJ4sbRRaBk4SNaDQw6q+yyA4x0Paxo1HWfKOnBOIGXtnxODNevkXFFbrh
L4KcLuUlX2SYtKzyWCB89R+jWPxOWN2B7SIjOzMymKAWAMBzX/QcdVNpWstJqd+M
bTm76deoUbjKtfXIKRsdcBqzg3ErhATeorp5aokZiZnbqbfZP7HV/FgU6EEzn944
p3Nh0XPIQz249Su36PDRu1qBieDEBW7H308E4g8KuOPxvhWKPnxyQ3GzR1+dsbEp
W97F2kFtxlM7Jy9nLVT0VuYIYQD7gRoSMKq0ibvom/Qc629ni/5NwgLKUXFHfD+0
uMGRPSuiUumeBuBDX7s0jsjynrF2i7WUbxpaUe57ZpywoKqiVGkA/IMPBWzOBcGs
L8VK5yK697eKt3qT8enCncwrefufMlDssRnUdut4DQBKT+/bGVapPnlqEXR9QKt8
fpTmg62DsPO6LaGK9p1YzkK0wMvjrqTOYCZ7UQNg87ALOsYwaYqgZ7BO7OxS2JOg
Uhb8zPizKYhCdzHFuWDjMq+WrI8zXVV1y2/yhx+5PvN9iiEf4e9lhNtaDb6iE7Nk
OZg1Y3N0DoYIplNKJWoEoZ9sccLX3iADEvVljyOYJ7WEk+Is5/QigjzuxZrwk8CV
h1S3+I21jNev9QUVLTwF6l+jHjyq3zR9ypkHN2wUD0PY6MC2F2Bb1f96pMVA+WtT
5RauFfz1jz9TQc94Ra4VlOScaKB0cRxLm+y4xbR5vEPP5O6H463Ste/P7iicTxCO
W43VhlDUZA2OVnldXcHpOQx0TdTsdHnBq5tbUKs0XRhUXDSs7GJUymzYaBOPmktQ
NeskSuyf7V2WGtKhid7OmC7kRcQ9sNhX1UGDHuuZFCHmZdMVqqwd80ckS+Hw/wxW
MF67ukoJl21sfr8ZKQVtjVknfSYbpWimgN/DQ7H2NO3OcChZOeNxpXi2M4KGsygh
CKTmAg4NnG08QmLJ4CFyAHgFhpWLQW9dcui2XR4TQOhdqHnZBVygB0RdF35nPJNi
nkVKB0KEstzKPZu7cChaSFMJE7ArjKFmA/p+JLEUvTVEBg8bKMykkpKWfrbnbvlM
N08n63NgMAT8pp3q1KyfI/z/lcuhBcq7YHSc9072Ia1rTo3+F/JgGD4eg0WUi+yK
mifXCt9lKlJjqkTzOovSZ1TajV6Du1G6Zjfr75RAgyZa2Jd2B4aXs89wCqcmSrKN
PzwkK9FI30u6KX9j/Z4eqTWkSrPHxMdC03VNG69Ev5FEK6xlZPEqGuULrUF9Rb8T
qUtsr9Ns/sZ4E4g0RmxIYAXcH5114A+5u3hRwFD//CxJmM/bMOFMubi/d2U16m4X
q8yCpj7qNBA+UupZnL/KUXFyo2MiQ+2UtnQsoyEBXIRtOHzQRR9l84+MBzqF8Ak2
/kxMOgcjGYP9Bgz2uYjRbYyi/g+pWdA9nV1Fqt0i+ZGfhi/b40ejr6JK/hCixGP/
eKRiCq4uc66we/JL8iJ67gPBgy3dmZANl2xnlxzG6Z6rTHlK+aFXR+2ailWg1wrQ
yrLLNHcnXF32tMnd9qILYdB8H0BLzEEX0nB0gZfwhiE6R9sS9Su8B9YHyMevQT0d
RMDSvnPDwuuTKdDXlR1Lv8uHniHIIhuNSUK8Djxul/n7hRYR0ET6OZZ5qJHwBn07
Yz1QdR1t0Aigjx7I5OL/5IoQkze2cnyx6SSwsCu6MoAV/i1AeijkRADM6OcmtodP
Yf+jSOWoZGh5ld7oXhtfelVp4EhbPa2aBK3RrJdmpWCkd17xKtPvbCIPZ/zYsT7S
czPtAM75Ekd5F3QCaP5OTHsVQv5HGv7CQEs41+KcmP3pTU3Ll1K+mcT9iXUGgkNp
qt93aF+wDtOgU/UczTgv9ldjwyBQUV8gZhPfk364XP6IW2Jd5TEy7Kmh54O99JKs
TppwlpEtTVe19UKNDCl4eKqA4qynvUKiSS5rPNpgn5AXgUgDltjU1UjGLRxWDZm1
NBfZeiPR0PJPjtlctMeUx2I9EeNwPoDGpnMOE53NWO7OqWKsBm1QcJ1XNpcy5eKc
oNeFYvVbc8nd3xgu5EsfCFshpRneLUsP41N4ifmqSs0KAZ9kUL+g/LOu/xVGm0X+
ph6EJPbW3vIUyfaUE2Y5X9xgxdQlFKW9zWx3kC0OW/lwBlWp06tcxpHYAt7r6VRI
AfUJ6iMnp0iC9Uv6OPX6nvd1tp216ZQCNOST+CheMkp94m4FhcSOKT/fiaJnx2Qv
dIC2EiPEDz1+SzFKnJYHIxo0X/g3klNMDVIynsZQa/yd7ym8k+Dnju6E43NS4UwN
IoJfZTYNjjDx8KMysvNFprHMwHltEaXCj11Ehgfrtv70UBF30saiSSmTNoKqjyh8
F5H+K/w8Tlxc36RLnFHDKDu8pgTnXRKbdCFbCHHIEJ71h1PkGhFdrqI6jg/Xdhfa
zF0KJVLgnkzz6/wsvEQEqZewEM6DrnsaJY+SlgpPjyUFn+RgIhEp8LdYFo26s2HC
tteNcKWie8oa+u5gzX1Hm37P5BpuoV07BezfgbIeQPsN7x3vxafvpvRLpzlb/Azs
05oKsASoN4AbPy1TlDSwxiWKuZnEMN5qSMZnaR0fHQV+oQOhR+LQ+2JRELekdOlW
RI+6VJ4qLufpweW7HIHNDH7ck+5mfFPJZ3Y2Qarn7DasIacBpIemOgUifCIpEDhh
e/NEDBAWUNUqlghvMrlbmIOe9out/sQBj+vVAQhKw14bQhRfAdTgAHTUMcnDlS6j
zN0Eu6LdexKkGINB/dlRt06m6J8pX+16PKnlHi95jZi0quiU1fn60PipwLQQMSRy
y6FgvIyhKcdf9bwfE2UUa5qqJuXeDiXoLsVwdVwZxlbJZAGcWtq3EMZM/zyYRnXx
IhdTaIywCkn4mCQRYH6HX2gZ9tJVtuBET7PlObD/yajjap2z1rJVFy4t30U5IXLp
gHgPMdIO7XVerf2lIfoM/nfY8F/gNTBpKRfSzeGw0lgp5LGt/aT1pix1d3uHGst/
MLwyd+C3VBoUSsQZhJ8WaPsabRV4M1NVOxDQffv+LmYyXr15IvMBvWya0HILl08g
vE2ypZIxTKdXkWIJQ72tx8xIycAznDAHusKYi1gyfCLBxFFPo3m1cqRyjG2bMmTB
7/7tE2veF1gwbFmQP9uJhnzdCM7Y3wdPXMLwcqWZZge4nfoHhCPC5a7RPYoszmi2
2AlNECxceMRGUYdf5hBYOw92SASeAkkg9gAWpNlF67xjpgHO44bSyw0CqQ80IRrK
5H+3Wp56Pf1WdRGhfD2oUZXh22yEyJGHw9zK0R9Wv1eGJRbP2ScXeRaG+bS3cI8c
gIcKnufI9tudB5hMEXIF8KP2X02GQu27dk2H2SwNMHYgLlDg4jKFUK6vWqDpWR1f
Wj95IWjXDsCnGLUsnPJsXO9dbmByzWWq849jAkwXUnOwjrkzVh2ilgI6Hi6PY4S5
zM6dy0b0M/nacJL4U/80MEt9cWbsw7vRkOLTU36hB0LIS9tEklb3vYgn5vKzfa8j
WyXwqjhpK1DUhJdIOX+0iop5yQ/y5pLSZz9HNYpV914SZK1KYnkpDAqrTxKhdqUi
r6jUuIoCdRxJU+O+tvLqfBKzGhmqgXKoUgiS9tf8+iKmnZg0QbwOqxN+kgZLS1Z2
d6IVhyQVZsMXsnrM+N2kWf5hTkQ+1fIf4w7uETPShNoMBbD4wUSTRCHpeKY/bJ/X
u4MTMTpdKIiJWw5+qW+cyHcDwkT8ovjmUgsvmtluLuQeVAe6jxeJNdBttWRF7bTE
r4+0vIkM5f3JOp9BSSJZyNFvAnuAaKW0use9h6eJl73HO2wN4sdKf+MoNmqJpp83
Sr+JhwxhWD8OKfh6gF+tmLjYXWPBSGaxXo9q2A5n79+/T6izvLRcX75ks/nePCfc
mH1I73T+g+HupTwpKDhmuRsJBX88xNVi1PL+Qm5HDgYUUpNOn8K8PRT09Y+Hov41
ChD9lwiUnMWJzSlJVSsZ+RxK1qrKOh4ELCecTZGu2760kjqF/zSoxqaK9UQhWxQ0
/6C75+I+M2m2eMmrVjwdq6pnwBRrjJhn7gVp9to81Fakjx7PDXej6Rx6xn8Wv92a
kpb9eh2D56Fwv78HFzMHzZ03mW6/sibDzQy+TKifxEKSJWBODqGcDMI03g/yxnN+
FcFQqv/lwXrueqb2aVnUAl0VCaJ7cHBruR6ya3VeSF61ZzmcF9io/iE0FtwPZmrA
F0Z8eNnJPPrChTf5jnb5xKyx3vXc9eLVnUgPxqY8mN/zSsuNQQYX/Y7Ztix0ddmX
KMhLY6w2yQj7ApNtePUFsaYt3Iaej2sZwjH79dlxl4Njq03YU4B/90RDQoveF9aF
lPebZwdYM4gdlBWagFMu0l3HpqARSX0CDajLHK2aW2Tu1IuyzJLpu45CJxKDBFwh
fyTzFl4q5GeQLDLQBWJ9U2nwgDdE3TcW1a50iQ9v6Oa89gWsBi0eij4UuCUEm4d6
46cQZzIGI9JcrfkycphwKN9sVQ+pb4+foRDP1UTuzmmJsRlVoRP1gzy9G8zQt2cL
pDKc/ICu0y1y++4+ZcXL+oOTow5iTvpLMgizHM5e6RTp7/GJcAG2YBDhG2ftzJO2
o45xoz4tLr/2LWtHT9bi8AicpLUI1MgKQ2FGw4VqSNE53ji1c0eQPkWlO+rgUa2M
6HZEcn0O5SJrsTbMcAAXs2ebtlZeCJyc/wZFz9AW/s94wDiUZbgzKsk1h0pXV8bl
DIEA816a15zsy85zmyO+ZbezTRX5dF+A4JqT80fkd7jahfckOfoNcKwrVLUSOh6A
XuGefdzyumqBaitgBMeknW2ZvoZB3U5eta86FMpZ156qGaQlxd72ZfWkP0cZaSx9
layH4pWLmxttPsZ4BeeOQ/kmXDmca9h6gYlzbyknf4IRpj7GsSQ2dlQRlx60fRxs
qs1CF8moJC+OCBDisWiPdORGHxSuA0vOHgJEKmXe4eq2TWxTOSZvlRNweVKcoPJq
VOWt01OT4r+UIlX4P9+YSiut6GncYiW8S5KqbqLDlZSXPbOsvCliJG4Iuaf+7Tbo
D29pa/IQ3OcGNF+YbG1jBbsL/vanbHkp/HZseSnSGi9I4+I9N05bJzRj/CPacMA8
00cjjnU7Z7kkvLPC83OlKHFu5vuNb1PNDhPfD6BLED2nK2UQ83MI6szlcYo6fcqO
Qx/3imFlK43ZHGLImkza1q1v228t5wvO7xCGNbdGrsEQCmRW/lMYR4/p0iNAuVVM
+hjLztN1jf4bUwIBy5WqnLNNp6Q91L3/7U+EWiK08vPhcRH8dfGyDpTQ+x9tEFB2
CCuSAb39511Lw2M+Rn/DvRqUdeA+tbwOZsyLJ/TwCyT7wm6JqkIo8thEEy/+6RLW
OMfyiOJ5wArnYC05qxKcEgP1pRRVWjrMGZ72Yf+jdsVu+R6CxId9odoK5IoQ0aKA
en//6+/wrm6s0sqzwQ9AJuTfIqr9/yZ/jVGgjNJY7QJ3IkLkOxZQ1omoKtvOoDTr
MEGeNzK7huXMv98jIybLtHp3eeK+W7tmKMzqjOTeGtwfIglLWuW6Yv6DRIJto18A
6WyDQU/Ag/zEyg2bp2H3AvFeETOBQ4wxjoaVe+To1u8RJu6F2XcnRT43w9eQG/oh
CPUAtfZmIuzmQtNPBtmMURXriAyITXTqVEq931H+3RcaqkUUBopVyIH/A2VU79cm
45FPXYOT/dx47SpTcMr43hT3Miu6iccG6oYlO5Y7azwyEPvnES2asRriX69YFDRo
mXJU2dfojBTwXer4b6FYPt1MwgoTDUKmW9Yk2COzUw6O9dsDs7edsGNFra4Ej2+1
y/zlxzT8g5D17WhkVSs+Esz/mSm6MXd+xVjn1H5p1nkPoAkbxZEudMklIDq252y4
Om3mdB5z23M02v1s7YVIjclpJmmIvbUKmBo7VXpPPi2XuTRn/C26YNCWMKfc3EiD
sfNgmRAoIJw//uaOU6WFxQGkOLLqVb+tVfcdnfU7VEF7Afiz0vOySreCIO22b8xN
gRvBi7ZiHyaTjmpQ6atg0/1GxDMrhaOotaerVta1K8NSUKMa9LbeJMwuUsbMIvKI
1Rm3j3F2kdbuQGl14vs8QD96k+KrKYXP6Q5hQRi9dw5RGJ8PSPpSIYH5HfFkTSXH
0Q5ZjonQmsj2lTJvqAE7HRwe4GPDm5ziGHg4ot+5I+x02Vr0H4NpfpbI4+6v7u6I
MRHP73mCvwg6qPkoi8E+noCRtJjFhFhbL8wp1wheD8Ya8hrcbGSDKILm1V8en6HN
NuSaXGuAdP57tZjOgsg6x7n5VV8OC3PEostvqXtoDXzc30AG6sehY8/E/S88mhr/
t8dB07hH8VyHlE7psW9/eIM/4HwpfKPUFkDB5NTEcW7wBMu+gldUZhVY/XpfgkT7
CEAmEQqysXQSkwla/3lMfkRYIwN19b92AyqW++JXBnuJaRsK2cKvvNmKed1lDisG
8oR0LXgBBodRS5tpH1aiG2eEP2NaVN8BbrCDDMC353C+wjpnWtjKC4gJtsz8dMm2
FxS1b5yREI/XYH2H/R9twHe6UEUhkRcQ+Mq71Djr9HYH/UNcLlG03Uc86kzUSLlH
eP4WssWvieZppmNSSVg0EKBVMxHfT8RH8Twga7DNEzLRDlUGsVTbuAe3v/8tEFht
sZugbgzGqP2KmrsoPWOj8o7Zr8ja/tmX9WJu12dAgIh680j3XnF0SMfUEXO38Jsn
P9/dZdNhOEnmfRsXudaxkr/1TcGj8eCaW5evZjgjH8baAMB9DFvA7li7PyGN+yr/
K4ZsA4fiBNUFOOy87GJZx9i64QlsidswJ+gqdYeCxqm1SoDhdIU9+7+TmxgIcs5S
mZ02J1dypE4I0RQIPZOvdMI2GAKSnhh9n9OyWTi7Yi3JDnPE4RsKZ3U5NoZMlt3C
RSvrk0zQKQq3367Sn1OsEsW9wMWPXdEus+Eq9a46f8RrGm6WZnjKzSUkownPV94S
J4qYxMl6Vw3YfC9kYmxybw4lefQtcqQ/mG6ixmcc4uLr1uo34PL7qUWsTKffvmDC
78V87nRYPZChX6QlKtghoSwN2b5gFgw+R1V6ykb3wxbvrd2FOsa7HFXVt4bWSlYf
8WWoKtP5r7p+m20ebRZFvTDXDCrJ7+JrS9eLREky+OOYI4Qy2W0oom3H4393S9xO
66ILvHXlrMJ+CntEKUmek277ISBjLfy2EAJAEG/kIGymKpolwcPmLeldUefWoy6l
tnJgEoTUd6GP9DmGubjk9f6HMvfXgELH3hqzXKyKxoOyi2msEK2+uLVlS40sLh/s
gvo724x5breEoc4hjYVF3qLKc9ZH4Ir0tvgZMRb3S6c3ZQtd+gdbnBrI5MsQCr2I
NQimf7R3xQb1/cluHU+Mvxw6OmLuv3KtFs3dDlJufBDktlbSl09+MxejJsJxKpE7
QA7jBVh0gVRYK2ebzhYYyFyPibYskde/9CmSU4KQ417tues8I7naZUCBl7yd5SsO
Q0bXf1ODUineuKlVE8OixxcIkbZOusy1W+7zlRBJM3AUjOnmtta0ZWyzEMRRDkeX
uYjc9LGu0lsmC40pXBMb2y21EVsCRgeUBE9iP/egfWWZ+5JuW5RLNyQdiO/pRhl8
dHg5FdeA14L/cqldrYlxyl5b6XZoBf8U0OlWWaIEFu7A9Wz7rNDHAhVXjicvfdby
boAT/s9NdjG9vzNQWu2BW6UC+jV1jhR6oZLW4wNg1yrRU8uIwAuZHjoizNjIlOl9
BsAmekIyseKXGHT1qcmsMaOkkY5GCToXUXrRNuZZc3+x/Xbt0S7k2pIQmPj0vajW
9df70B1ivJZmjT7jvT3B60F7+VpxCgNjqaZRepYk2uc/upF4poW0Wbisu6QK/aI1
l/e0jzfthQDqB1MM6vYd+77XRyjasZxwxUwnn/fq3TaaN5sfmDaS45juSPwpa9cw
IIWeAQiXmewPf2wbJd73e/Ub+lKAEcLeq3QYnuDRiHMWc91pQr5IBVeBg2FAFb0u
SPVCzcYNeJST52WOF4uuwxqNRYbGmhFKBHZfjIt/wtcMSQFMSYO755M/lvV4iKVE
Bp0LQkkAaYn9RHFNSmf8gjSN1BWcqvKwIAKqYPcwf6hckPKjKSvWiFuqiHHWxkb0
BL43zHwj5bFfLCE+S4vX2afsoqEHGeupQSV2B+HMqyCSfziI1871WNGGG7imsYLN
pyN3xFh2FXco5qK6SOP7fQRBwL+VBX4z5iGo2W3zvXFD8sPr2JGvz5lKPLRth8XS
DRr/UBwyxZiN1V5IQ4nRLy7RVQAp4BUFAU265Huwj3qR1fggXg638yIv4R7InHSX
zrTzUj9lYKNXmUhRNNnwLKhxupzsH2uUkhkSAMlRPKR0999TksSyohXheS4iRqY9
lcqoKtgwjTxubMV5Kwvf0r0ujozxEhBZspYHi7A3BvqbUTf2kbu+VQeDYDoW0veA
Hzjciaujkn31T9iTp3097h7uzCrt8urY0bxWLTxapBVr9GrsmgM2L44CtC7bwZZy
RY/c4wKD8uGxuv+ls6asDeuWxs5HHUrjHtyC0BjL6RRXSrpG6yakl6+H1mt9Jg/g
XEJpPJgR0Kz2lvpiv2gWj8Gz1oNGaaQfeJ742kq1OwCwRfImQM9gSnNSpgaeHmSi
20J+GR71o1RbFL1/HemsqY2MiK+LSIbyNckZ6QCxpngTMOVLvEXDj94U1LliptJn
Mns6l54wDcz5VB00C4f3JR8wk0HHIkawbmRZc3ROnQ8M8aKZiP+gEtfKOrb49xQz
dFo3cAC1e3wo9toLAQ5gUu/2SUEVMP/zMu8d8FGH3sHX1rY/kOLLMX9GRO/wj/qF
7Vkjer0iAMaS6QCXI9VkCEKsBgY+e2Aw6sRocluAteG/nPOtlKaGDN3ewcXsGwKQ
tkUU5t2+QEyQAd27JISAMVR7Nb9anESvmBdoy1T8Wzfaq1Uci5+l3KWdqn1fOZI6
PiNi+a8jO92vrp5s4eb002l8n2pCLZmHBylpf15Jzab5a7iuPe5E6kV55c1Dhy/I
x7hYQAKnqoGnQDtOF/mFLH8CLqXiFvDdYlK8SnU1PZTUhWr1Cryi92EP2OtdQMBl
gBQYLckOCuXiz9EDeZVmUKeBgEM6an4qFWIMVe/EnttdjuecBHq0sQFVL8mNj3Ie
RSvPzps4pOw4fsakZOg4o8ZN3PyjKSy/neuvahFEmYatSJm9s0NJPgxTMrQOt0+p
4jolydjklMjK61fh4FnStoN1XYqCAYWEVzHOwrPZcD98Iqg80qZYLo+ezvYmZ8lg
xKhPMn3bg0bwai5cNGaHvuNcssQzmciIB1/8BdrKab8/lpZMgLzyb52JsQXI92V+
wHp0FtdMEN1C3YCIaSG0Gtv+CVtJVpwZwEuEDqDB7z5ekpCUG1xIHmSGKY4br3Ef
RkXRTF0/O0czupA4mTNmpxUjAc/PimWvetJ3fgYJ0usWHgjZojC7BQFZPNjANCNF
GJ1nGvivLz0HxbBCr7kU03++yb2d7Df8rH4wn0W1j0HM3c183Ch94h9Ow8HPgpzF
T4Ie1W1FHuiJuqAAcz41qhDqnfxGICDEpPqp2o0BE6dJwxM9Tv2t9Bu5E4pddydC
0BoC3ojwt0+eDp48KwIwYrfCpf3SAoYL6CKZpM7+06Y2EI4krJzJtELCWi1YneBF
qM3+KNeTEuIYMfwq8oMXaB5xJhh2e7/Tl3oTwbYsqMAsDLYsfL1IkD9w7ASVukZ0
wv2wP1ad68CIKFkKfdiTJ0CUYRSQinCkPHFio49Cnpb45uoObQYXqKk1WgZ9xfT9
UVDUVlqM8LNNRwx9OuCQGpd5zAG62oHwG8k3qiJF/sWnqYeJ1Vv8F6Vaslt5hQx7
DVNOegsCdwAvfaoSemfL4EKkHueYNYzvukSCV7zKIkjO5xNiELsQGx6JiI+jPV0Q
dW0XNqA2BEqE478qR1TN0A2I85jJeQVhjC6na/xP9Lso50rqa3SE8spk0bdRwkiR
9JVP87txot1FywyUe3JUkezORxCPbAsRTWskZvliLh+Mtn37TbFN7P/jdbgs9T6E
S0nODHcD2um0LIA6uxhHAJBRJ3IDX4MKti9irS9995nE4uW9miQqOawQap8pj9+x
UkXb8Ns4ns/lzx19BWJ2GWZXY+X/U+PBWb57+/ff0i35YcXbTGBYoBmferBwsHO7
9kcTadmXqsELBTCUZF//XdJBkaaVrxIENSp/MXJH8X1vq3hrn+93n6n5evQ2vO3f
ol1y1gVdC2Ozo5+RrocjNNwi2Tc8trmayV23CLDoVg1bf/I8K3TkQuQpDWLFBiTc
GIMEvNHx1a4d+o93RF53SSFn95Z1pIHOwGary0Xn5TPi4ehq7sdOofOQXs7rhPKt
aKzIGYbUkBV5IhfS7lYM6Cn5TobZ77TGnGL/i6n4VcV7zBFYhEYS5rqE5UZmXGzL
lNQWcY3FDCdGR+SXJ5PqerlYRP3SBHO76oloN0WgNYXQhn4k6t99I6vjlEAH31sC
zAQsIp4YWTDMtaYPH4r3PHpsdW+Br1+yeUbEkGS2JhC76qDxbLScliKEeGWC2emQ
ouHMw71xzN8AzWUHnMp0cZHwORV3ykacUwi/sFb6LdLaQUyhTcxfE4m3fZrdBKdZ
8oGk59cBGq9/SHJM1gGLjWS6UOcdz0k5T9aRRJNNfJsVioqmW/pAejJRAjevvifo
k5reMfOKDo5UvJ5w317s5T5FIVQy7AdULObVL50LZ1mCetePdw+U9Eb6juGDw39/
YOluUUDj8Q33HmO1PFNd9QmzbBvBvNy4sFMccTc5fO7K9f8F8QeRgsgE4L7LOfsd
hJb9D67rxLXE6YtsMQoHiWmsDV7kuqPrmfNXC9uFq+FYvJqPzvR3whDxM8WB/TtZ
MSkQHvL4Nz2hEZ1bwweznfiROYPm/v7PiZU8uvddd0yniW+Lx0WX98xr90DVWl4+
TR0rjOHoUV/MYgEo03ljUVgrSwDWRGbgaJgpiRyXT/L/POCUqa3C2/Bl2YGCw04v
eOmW1/4WC7Ax0DokkTpm+62OST6Nav8M0Hv/YHVl2Vjdwek+jdTTmDoKItGwzUlv
TLTvuj6TX+JQwHVS0S1ANUGURz2oRVgOJMLYpWw4P15eZwfJZBnctXTJRg+ngu2X
5Y4rdWwMfu/b+1BehpBD4yJeXIVVsoUrUvTLcDWYrqPsSNzOpENtZhvwlkx7VfuM
GoEEPHY5P5f3V5aQfoJVyL7aFtVAi+mio1kd8iZM2w6il5v/pwMvIxcFA+kRpI5v
lXTHLORZoICdqRkEjwQKZroFdIWpQ5fziYFY9vYYIpbGJxGysyRvH4ZcjNqzXTFQ
9bffPEnpx1IvtJsx8V6zQfKscqWceMpK+8NPShH3BtMPQnvTBlV41UU+/r6aPwGz
nBzIJQn9DYmGXumaQ+U/BK8+3zoBQzlzo3CYkwp6W/ATVjcT+1gF9G5DSnLrjAWf
cZn5sgzE09Gfl2/eVvQU6zV5mtDh+ylvqpPGf7nWFgwmqm5ks7oBk9vmlfp2BtSI
9/m9PyZ65quwBINuS/6RkIYtyrCPWDh5MCL/FSVApJbTBtPFljLmb/Pdv5AY7tMj
Ck0NJURJBOEtTvAtRHJZkUyV7jOGndRC6dHAQXrYSqzL0U3otJQtto7G5SFaELGc
3+I91i8AmoluLxwuUPVv6Wgi4uiFeQVwrZdejDyszOCbfdSxzq+zq2ib4K1w7HYa
Gc2fl5HlhKmCjlYfUtMCq30UNTFmpboHy6zmTeALWmAVW2YBfBxVXJT4RnxmXeHc
F373/zwji9ffFAC/7ZydG72mLYLFjUdP/v1wkBIAq4TZhipZTXrzZcCd9CpQ/icJ
ApjEzwbaJxOTGpqx3J+3mFXWE0oGRdR4mHgSWTqgposRxq5bLr9g7DfDVBNQzh6y
EHepaV6uJ2qBjL9F8lEOQQVr57PNLcK2f9RhlwQ2bx85vk1leyT2hR6KPfovGvAi
yHBQWiAl8UM+DvuDYnSt1NKFFi6pGf3w6UGywdlM3TgVBdlDw0mb9U3OVU+HVNRo
eLEL4lDxTfEZzKPJCxYLYb5YnQL07H7B1fqbWI69S84fEPKMbi/jwEHmSoTDeqbM
kzymJaDsqi8YfOas0draK95AQMxWzInA/5sofUJmZqwb3MHNkdzSYxlj7fdKAAd+
3kMFi/Ud3kRFe/S/n1qT7EvXBOSD3CEkPd7QpZixWYsOG9S0ih2zlnEiluCqygzT
hNDfGGR2jsF6iXvaivAXdqbniBJLhsrWtpvCL0iuNJcYM92WjAgTGVT8r/qZSVws
99yXB3j2/Iuq/N/2jsoeQzcz1zgm0ZUHKvy7SoV/VI5Y/IpqcKjPh73Uaqc/y4e0
MH6WNGl+BJXS9N3j9Fpmthehm/LivwctX0MKjicUFMA13jN9iL6m8FU/gqedsvjr
7UiQz5D1nQR4ORIaD5gSQAWVvtvjiWB9zf1I0s7/USCUkukkZ0ZB5LireTiw2fTv
sGojYf8m2DibYIODTxNR3RO/cID3wkEJwAoN3/rKjCr768t/srrVOFQz8czOWn5y
caaBHVbT9t5H9VpUpig7Y7ds92/a1VoBhJwOuMuCJPSNCJ/PY/KC0Yj8G1nSUqAC
gob5E18OKEgtvEIIxO8Eo9xNFH3W6YQbBXiRF7mAEWIGkpCMLCp4XOWdlTv6gudE
YgsIu/WxODrgltwYSqjRnsVtzrOrk6o9HQOr/rjv5TSVIN0IkA+EXsaH8nmP6tZR
A+cFSuZc8boWRkiNdCkrQGEhteIyiBx1S2YZQM3uLwN5/w9mI7Ljn7iDeMp1ambL
fohA7wxKT5YSMuX3PS2VKTVWFqqeSO5Cw8KclRXuLayjCNHlhGCYf/wCHGIuF3xN
rl/X6jivXmeiC4Yz+7S2OE+gl3IbFsBhp/Tr30WSL+x1e6w6gEfMxr3A0OLFCDXt
WKh4Gb4TEKttnqfjQ4sfs/RdfygajA/sdr06ND2Ohaw=
`protect end_protected
